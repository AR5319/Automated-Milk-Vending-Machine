PK   ��X�ji՗6  ��    cirkitFile.json�}[o�Ʊ�_1�_�A�/��$�\�F|��`�����u���x�ﻚ���C6�8U�dDZ@�ͯ?�����]��z(���������ۇϷ�wW�����|h~)��*��>���<�������Շ�ߋ�_?�E�ЖMu��X�[�m�|��1����B��!�h��7��������?��k�obc�`�,T�ua`T��E,�ΊRu^T7��z�^kTU5�/��e,tQU�(��ZV�+�&½?^_N\f�7�R�q�pm�&��(;���>��x#J�y�x��JWuUT�S�	MS��n
[���^U2��u]yT,*�A`��E�X8��4U��S�H�](�]YTmh�E�mTeE�^]k�\t��D���V������躓�(�����i��� n�A�h2*��1��|���o\���dE(m�DW�RjinTF�p7+��QG�Y
sM��r�#�ZK�V*��qdTq����&�9P�M$s�"�L"�S	X0Lh�Mҧ42��Ojd`a�,�"�k2�͔t�I� t�I� t�I� t�I� �n;�"��d� C8@���n;���n;���n;���n;���n;���n;���n;� Jmt�*[tmYF�X��m
��Ayن��~��� ���(H2@��˪kʢ.M� Z��ԝ(B� �l�����dBjm
U��F�5EEYXe��/ �/>5��m��[�c]�X���u��5|���]״�/\ո����m��R����.�p����G�����h��@E�h���HT���$*��r�aq9Ɂ�����)�0c�����U-0�`	cW��m�1����6-A��|D�X^���B,/�`YЭ����N/�a`Y�-����V/�a`Y�B|���}(�ۏ�қO�ˇ��_��Ϝpw�߈p����eo�Wv�Wv��$/;�\ye�xe��N���Wv�Wv��$/;�xegxe��N��Wv�Wv��$/;��xe�xe��N򲃈�Wv�Wv��$/;��yexe��N��Wv�Wv��$/����3G��$3��v�,?��;�`�/$s�!�#^~��_Z/b�s���O2�K+]��c�4x�If~i��Y~��/?��/�.2ˏ9���'����0f�1G��$3����,?�ȃ��d�R���}����R2!�3s���O2�Ki���c�?x�If~)��Y~�;�[��b�?s���O2�KI���c�?x�If~)ݗY~��/?��/%*3ˏ9���'���kf�1���$3���,?�����d��ڙ����g�=�O�RV��m!}�L(�X6E�t�DW�����d�ˠ��׮0]e�ة�0UhE�T�	�F���^�u6�ӵ����C�붭!J[��h躒E)t(�3�7e���)]���u�i��ڗ�!�;q@Q�������<s��"�|�{��vKynl�zv��M��'uM!�I�+o?��_;���4�|���a6��^{�<�7*7��>��^{�if���O�aY{?Que���A1�D��|=��~��O�X^{?q��|%��~��N��]{?QuUNuq�
	���#�3Y��7�!��1���%��2�p���s�2R�tMs�h}�c+�ǉ`_)�I�%瓠NV����t��ǖ��(3�c�$=6��ux(�m���=��>7�O�s���F!���F�AJ{���F��s���=wn�y��6z��L�ύ������r&���a��5QOs�y��+v��1�ne�9�p��:�n�ǂ�5O�1lI�Z�d.i{
�H;����)]�^���<u��B�ھ�u��U{'���$�����
?�M'� QWT��Εz�މ�ba�w?q:_X���Oq+�����&�ʊ]���M�[s�?�=sJn����,rw�kd-�m�SdQ�m&F䁔��ѧa:�>9��L��4I�(������9�$�My�6��:�t��F���c��緹qg,�n�oءn�{P���������=�>�n�{O����R�3E�pC�b�)����ԉ0g#p��B�~�P��w��~�`[Ȅ��On�P����
����B:�~��-����-Һ�	5��IVK�ݳ����cf!���ߏ��z�T����x�@��y�oR���E�1��Mt���.���ƈ	�?Ο�P�?#&��� j�?#ã����<2b�� �0b��0b�K�0b��0b��g2�LHá�L���d3�\HÁ�L��l�4l����b L���d3�\HC�D&Nl6\�q.���"'6;���8�Pg�����瀳�q�fǹ����L���b��\HC�F&Nlv\��q.���#'6;���8	_�Hra�P�Ȧ4F�/�2"��Λ]|�DF�.�j"��&_C���y������輹��W�at���-�0b2��5��U���L$���3�LH�5���8��n.$�ʊJ�L���7jeE��9$z�Ev���2�i�EvT6��B�쨌r݂�:#�N�fGe��\��y$pzv0;*�\��:���#��3��Q��i�G	��5̎�(�-�N�A�H��bvTF�n�uZ)�G�g��2�u��*�<8=���Q�[p�V����Y�쨌r݂��$��M�5�����orm�v�@%?,�l7
����&�!�a9e�M�	ۙ�����&�ڄ�L�K~XN�n�m�v� &?,�l�	�6a;S,��S�ۄb���)���)�m±M������6!�&lg
p��r�v��l�3�9�a9w���6a;S���S���e���)���)ۍ�Ķ��&5�a9e�M\�	ۙb������&.ۄ�L�P~XN�n�m�v��(?,�l���6a;S`��S���e���)>��)�m�M��&���6q���R4�҉��%����0���A�ylUЫ��(��FԢ�G��\~Gؚ� �.j�P2��k��a�K&y�Q�	ŕJjJ����$��_WH%��P2_D�D�|�V똔7��Z��e�?�)��6���{_�IU_��Bh-�ￃ_�S�u)��6_ãŹo�����ܗ�kax�8�}�Z-���p��̺���f�b��Ц�0�����.���G��;�P��<^�x�� �3.5�|"�x��l)D�;E��l}Bx�F�2��bk.s�L�UNe|Gl�����V�I\Z�_�rV.��z�%�NRP�r��.�le&�֮[~G�"t˺�-(�l�u��4�F�\2g;�D9;`��-[Ll6.g]lU��h]am�!BK[�d�uϖM������r���˒1��!������U.`t�/�wv�F��Z���u�8`x��|T�.��s6�D���1Ź���κ�Eo��ri](ky�]�jy%[�j�k�V�Z6�ؒRgV���D��"O��W��B�`��a+/-s�VQZ�-���[�h��FѲu��*b@9�T�-\Ārvb1b@9;-a�1�����%��G �lв�B���<�{>>@�����N�JA0<J|>>@��a��<Z|>>@�Z^�FW	Z�A�Y��E�������>��ǖ���]����xL�>@�Z3#&��0ZFL@�a�,�����hY1�Ѳ0b�ea�4F�	h8����p-#&��a�<&��j�m6�-�7��0ZNl�[�o.��a�<���d3�\H��><��l�d3�\H��><���b��\H��><���o>�͎+6;΅�/��É͎+6;΅�/��É͎+6;΅�/��É͎+6;�@ZQЇ�����#& �ʊ�>,�Λ�}X�7�+
��0:orW�aat��(���輹]QЇ��yc���#&S�YCYSЇ�D�Ym>��f�+k
��pb3�\H�5�5}x8��o.$�ʚ�>3H}�Q���Pg
�p��q�)�Í�(�-���a���D0nTF�n�u���&��q�2�u�3}X$09	��Q�[p�)��"��)`ܨ�r݂�LA	LN �Fe��\g
��H`r�7*�\��:SЇE����Q�י�>,���ō�(�-������	��%rx|�mB�M���a���Fa�6q״D;,�l�	�6a;WЇ�S�ۄ_���+���)�mB�M���a���6a�&l�
���r�v�Pl�s}�a9e�M8�	۹�>찜��&$ۄ�\AvXN�n�m�v��;,���6q�&l�
���r�v��l�s}�a9e�і�6qٴD;,�l���6a;WЇ�S���e���+���)�m�M���a���6q�&l�
���r�v��l�s}�a9e�M\�	۹�>찜��&.C�}>�]Ї���^����}FA����}"tA:
���E���dr�W�d��W�d�|W�d��X���"b%J�+��ZǤ�<ڛK�_ã��$��0<�KU_ãù�����hq����0L6�G�s�t�����ܗ�kax�8�}�Z-�}�v���bͣŚɕ��bͣŚG�5�k-�<Z��j1������Q�rA�����.�CG9�]Ї�r^.؂>t��\�}�(<\�N�>t������4�.�CG9;	��0h���h���_Ї�G��G���>0<:|>���a�z<Z|>���a�����Q%�����*�}`x��|T�/�� ��J��btA:��x[Ї�r����||�-�CG9�]Ї�r�������A�.�CG9;1���Q�NK�>t�������1)/�����}`x�||�/�� ã���|A�ǣ���|A->��0��h��� _Ї�X������Ǜ������m��__�r��~�������������i�>|��s�|8bM�B����焀�l"��P��U�Dn�P��T��n�g�F.y�v�(]k�����)"��6d&�mZי���d)Jג"pM{lIQ4ES�L�wd�\�gd2$AञI�:�5r��2�q� P��^��W}ri_�w�=W$�T�ҳC�An�6�D�sdf
e<�3.��@��2/�&����Aڲ%�L��D�L����'ѬezG�\m�9.�j�Α�L='�s�ѓ#�g�����O.�����yrl�����s(��T&&�����6D��Dф6o`�K�w���[���](��� ���m:G�n�9r�3���F��|��l�@!��Rפ�� G~ct�m��8�H�%��H�k��d!��Ll��R!�mi�0[h9v�fs��{�=5.���ǐs�q<���ÒsP�U�^�sy��/ %h�b��0�:�/��@�Y�C��8�g�aڠg�a�����C����[x�w��~�����w�o+��g��(���3���t���E/�Ag@Ά`�@L�``@̍``@L��3 gJ0P�&L�)�&	�D�� 5�b��%S��Ĝ�W��� ����'Z�-C��$�i��IϾX��I�^ �a�$�d,2x���1IL�Xd�"y,Ƒ���)d�Ɩ���A�d�.7d��y\1TK�ⅲJX�kbrɢ^$��L�©'��LFʲ��Lbʖ��)[r���,{�/���`�_>E�����W�;t��������e@M�Y�c�|�Pe�M�s)���"�Wt(�^��8[z1�+�qJͼ"��\�HCˠ	��/���`@���HN��n�@g�m�a��e��q��/�"G��rT�9���O8����$�R�ܽW'qv��e2��U�V�^&�pq`�Dn!���QqKo?Kn�2�}�)���Kbx��r�=�����o���*_"�w3��_`p2�r{w���|l�><�~�u����͗����?i�	���G����ަ9Eۇ��1t74Rd�%JdA��Q�Dd�ez�����q�tI�!D�*�B��Y�!D�+�B��Y�!�p�,ը�1�pR-��u�敎!��r�<,l�.�C��Ry0�Q�`H�b8/�ʃ��JcJ�É�T�T1�S:��L����V9�U{��)C�>Sy0�S�`O�b8x�ʃ��*{J����T�T1��E�ǒ)D.�!�#t��d�#�"I-YE$)2��B �bX � C,��Hd��Pɂ��#Y�!�C}$2�r��^�>5��#��c��m�0�d�3�?��A]�ڱ<L�bԎ��`T�v,���cyL0������?��38�x���d��Y~�Y~��$3?p;�姘���O2���Y~�Y~��$3?p���g����O2� �Y~�Y~��$3?�������O2���Y~�Y~��$3?i������O2�`�Y~�Y~��$3��n��@sG �%7ô��-C�(�=�C$w "�#f������#C�h�����Q�#s$�;"af(��5>nrG%�%7ô>�-C�Ȅ���f����e��03��SF��#f���a�f�!w���Pr3L�x���q
3C��0erː;Naf(��Hn�o�p�)�;NQ�q
3C��0e�rː;Naf(���Ynr�)�%7Ô��-C�8����f����e��03��S�5���f���a��!w���P�c��N��#u�9=Y�g�9sY�h�9DYc�mu�����r��$�uu����(5�&���+��Jg�ȹ��̄���
;s����.w�n�2���I��ZU$��$�z- U}���Op�|pCQ�i
���� ��!�P�RN�B��/8G����k�z:�&t- ղN��\@U��w�k���f�R�L�GD)c�g���!�8<�w0���VR�XS�Xϸ���̡��C���4�F�/��ȲS�ȸ���;˧o��jRM�2�,�����ZP�7�|*��ȊX����d9!�쐥�&p�c�pv��E�&�"3h�eo�oYm;*pU��&Y}kB��&��b[	w�d��p��>2�|��\0����,6�����:t��X[�k�pxa�f"��c˛�9�wU���˙v�¢��#֋�Vu]>s-ތʓ�*�9� �6|)r�P�x)r�P�v&T��I8�K���px3�$�d��֊�%��+��8��"�.�Z��x��)&�ɞ�˭����ay�6��������B����a\����k�s�i�/Lm��f6�1����5da���p$��؊1XÅã�������ӣ}�PutiC@�ҥ5�����STC�����j�R��8�]Y���n�`�bw���j����>h�������&�ϩ&�����W)�M�J]�x}���y�	n�l��{��Jo2y&��8 ��ijH�7��U�&�o���s��.y���/��++�zO����Bn�'��ӿa��P�~�Q鎾�h?y�N�C�;t�C�;t��/©czL̆�H.�=���m���������q��������+<&�D�5���"@݀�F7`���z{=�X��h}:
o*xge)���:�h2m�IuQ�)[���� ��kA͝��աe���`�ve��j��LQ7]ӨNY�CK��+�8pƷF�2
WY;���l��6�*�Ih�UQu���f�U���1��6H�HxQu�qm�*B	d����L�C�X7������"x��nLc;�J�oY�6�N�тWd�N4ۀ5*�Wm'��@��S�pWji
� ���K��kSVE�d�,L ��rFk����{ X&Œ�Y��젓@��L�ξ�h}�J i�d5+'�����Mm\ T�}�B�J����@�-P�`>x��AKߩ����F�Y���':N�~U�u0��в�q�xJx%��u"u߀FU��^���a�t���.��+Ek�kbzqU�!0=f��1M�7{�'?iX�x��eR�Ɣ�̰!�F&;�\��(�`)�!2ΰ�6��JR�ʔ���ɕi���L�Xʻ��Ć��%g�xJ��ܛ
6�x='�H�C�c53�dΖ#��/gcg��L9���!�3��WH��S6cc|I�B�)+���CI�!�L߀!�A"D�3Pj�i,Q�2
���d�Rr8)���é�s362�r7%�������t�)�|�eȴ�)��t��T%�M�(�lM�0����M��<YR&֔�"�gZ�5%�w�,���)
i+cJ';��+YQR,(�(��	Jj�T����i"i7iJ'ge�Y4�}vJ
%�f"-�z��p�M�䂣�����7˪�������Շ�?��_%ѝ\��KrzI�/��%���������^��Kvz��/��%��䧗��R�^��KqrI�!��O��C�!���ȩD�A"r*y���Dd"�B��ȩT�A*r*y���E䢦rQ���\ԓ�L�rQS���\�T.� 5��:<��>�>���c�����h@��u�7o??��rt�3����Ѷ����M�;{�p�����Xx��_����M!���x� L6�	��J6�RE�
���V�E}4ֹ�,�P{c����)���c�x�����Ǵ!���O�>�jo�>O��Ow�?�l����p{�7`sW��~OW���^~��~�C�՗�[����?�������C�X�����_o?�Vۧ�=�����C�\}xI�6�\�}�����C����q�g��)��/��_�����'��Z��?�>�ރ@�/��~g��^����.���$�A����櫦V6bJ�a�	1�� �k���vR6WGo����y}u{����� T����=<��c9��ۇ�c�ˉ�W;s����ׇ�
t�L.�s�[cFw�������w�_���'�Wr�w
�U�������B�>���u��e�îPƘ�t�[�	;���Z�U�ղ�Emm�������5!���"TB��E��RPcX/����8^��;��t��G����<=�7�O��V��5�2`�,j-�"	���T�w(��ryP��E�5��>�_���������e�6�¤2�䥥?����������h�����*�#�0�&���epIp�k�<�-r���c-�/5(Q�l��Y�*�\�h��.�5�^6ǝ�N�4=#���(*�#=�~C4O�u��&�N$��2���k�- ��ǌ��6�
Ba�HB|x�"�7].u#QbD�/����O��H��2�k�AR�B��+��<����};wym�Co]�����D�x|J۽x��h���(������|x�ݾ�an�O���6��"���z獇qv���]? #���J�ث��]��R�6�\ѡ��;'�vj��x-�7�����KDm<����.ڡ��W�cx��L�`[�ǌ0t��H ���!>5%d8p�(p��>�������� \(1�݋�;i���H�T^�a��i��f�����ǻp����-H��r{��<�AY��*	�)8d� ��o�oΪۿ|w�#���P0��RLO�\8��v�5J����vRg�|���?0r���go�M��� �9�7ƥ�{0��	x�+;��҂"�g� ����HV�����}� �$�1��r�X������gzsx�qб�&�ð	E���6g���ah��!C�D��+�0B�dc����]ځ�����-�0�6����t��7��p����?���{��_�ϟ����ׯ���_PP��0Z�����Ou�x��kѩZ
�#!�+��CQ���]�X�k�t5��>�@����;i��?�pA��Vګ�_��s|E_�GWT�`R��:������f��l��GqOW�q3}ԏR�WD���:j� ퟮ��=n�f�t���i�8\�'��a��l�f��f�m�݌t����w���Rf//o����5���BbF���w���r���K6����w���fr���;�݋I�ϙVpp�SX4���6�� N�;�� ���8s�(���9���U���-��eѴ]W���!�qU'MS)��PC!�&�N�1���0(�0(�a��Y�-��d���q�<���Fa��X�.t�}��EY�}m�������@fz$����$����Vϵ��
��sQl�b����M��p8	��zE~�f�~���j$-�������S@�������>.����%�>]�}{	q�>�D�ˇɮ��{Gp��bt0D��d⯥Wi�CyG�́mk[i!\P��u�N7ܡ�n!N��g�O��.�*f{�N���d��ə��9\��ރv˧��p�	����>_Iފ��O�CB@-KOW<8l>��c���|���a���K^��i9b� ����}�oNe�:HZc�4�z�a�3d��$��
���Q؟��}�)$%8���Qap]A����Hv��L�qWpe�j/��*������]�58��Oe�u��f��&]�4w��^&�'�L-@AB<�/h<����H�.�z-����a�Dx=�e�ۤ����G]��颓a��hI��?�6aa!���y�����᫯���Y�ŞC�#��?=�p��}��ť�qG�W���O<��oo���}��ۧ����MU������/w��?��>=�9m������?��|�7��z��s�Z=u#�S�c����#փ��̺��{�����Yԧ�O�V�E�"Q�������s���S/�'L0�۴TJ�;o��
�&�A�(�2̅�x�1��La��/����O�����^
� ��^�ˍӯ���}x�ϗ��� �ۂ,�Je�ܹ�&J�6^6���C�����_������k�����U���isT� �W�A�k���6��`Ѥ��o2DQ����!�헟?�;����ӿ���O���9p��ׅM�HJA\�4�M�'ꬬ74>��������2:pfC������wB¤�����N��toht~���+�>>��Ƨ��9}Zew08���l��Sʝ��{��Y���oQ�B����G��}�*���f�U\�`����w٬sBS�6���X�� ���}��� �yl'��F�o`�L��R��uQ�������S��� 5��}��� �)GG�)`إ��]�q��>��U0[�kԾ����4��uk�`��"��>u�k�PQ�(�������t���}x���4�	��M�҆����O��(�5l��b�l�����z�/82����֋���;��J���CJݕ�MT]�744ߗm߇�Mm�N��fΘN��鬉]:�C�k)�C��MT%�746�Wl���ˎ��N�/����WCә]�"}T���mR�P������K�������/����q���4h��J���A�d܁���������V�黫�>L_xT؝�&T��k}�d�$6}u	s�6n�\L�R�0��UR�~x>ރ�_0�� ��풘
%��)���
�/���O�����8߷���?"�p4
�3)V���cr��.@�uY��6x:��ۇ���׿޶��������� "M����02D����~�0�����./�ڣ�w�"��k�P��+7 ��|�>�߂�*����?\����M������ߧ��/z:��f|�Pjq=�,} }t��s����
eO���W��b�舒AV	|:��u$�ꈺHGƧU�udtL2�����4�p�]�������~)�I3o2f���������p����	g4N��S�d�3^�Y��ܸ���H�ұ���f3�O���36O�;�ʆX��e#V���\tn��֑�V�$�Q6i�,�̛�it��Yޣv��3�2ƦI�X��)�fw�=�&���R��f*c����^����j��"i��%����-�������z�Dy�|t�Ldl��Drt��c˗mH�E�[V��QA��-ɫ <�V�a5�n�|��i�J���|󜓇f~��s���4Hԛ?i���/~Tc ���\6¥�Y�F� �'�k�e�����{q�,��mx�Ӳ��sI�eRyPɩ"�1�����e�e��A�gTd�,�\��\�gM���@�)�Ԝ*b�4$2+�eՏx�$cp�̸Y��pT&jM��R���Q��u�A��z'�z�ƪ�
v����zX\3n&��s>ȡ���f��flL���*�����х� 
�2Z��6�u֕5�Dې͐j$U���FG5�Qe��A)���ys�̮���*��h�7�T+��T*5�{���Oo���������]�j�����n�(h볂*QQBfol���R��0z\�nT����Tgw�)J�X�ꢍ�S�r�qPJ�Z�L�ܮ�x,�ݸ���W���R��Wt,�Zei�G[��f2�qTwM�q	�߱Z��Ŧ���U����O�Jg̐��������(�j�Tr�����k�Jp����k<�5\ij�o^_������O<W�^�l\��w�Tg79)J�뭫�v<O��c⺾���c4l����RG�W['�J��$J�j_W�J��N�,��(M�����2zU�-�ޡ_Au��y�C�Gs�U:�v�H�8��p\��mjU]yT,*��Wо.J���E-M�V���
�D��w��8ת��1�ڱ�aN���p���{P?�J)�튶%��������"
ۨʊm�����JT��)K�Z2ίh�pb���r���N�P��g7z(�ǻ>Ѧϩ�e��OZ�Ye���n�]�EUѵv�EWhȿk������ �7����L�}�T��2��~�j>�3z졡Z*�I}���e���Џk;%$�K!���SO\��߲^A�-
�h�z�qg���?}�Ȇ2��b������v)���i�Wc�F��C��UiE��
j\�tY���{�i�I*�aveU��Ǳ��$�/�J���/�Ϋ��eT%������/�^v��Td�y􊆙l�B*�w�*��I�LL�g�)�Nb�P��6���VpcӦ?.ANr�4VC���o��@���� ]����NÓD���o���V9���%6��Ix|�����j�,bYwV���b��V̆+��9V�M��Ā�ǅ�:���r�_aw:��<��`��^�ƝI\�J�J�q֨�j:_DS��4]TU�B��P����j��ύ�x�K��g�٤�:���,Z%�0��f���u�U/�(�u�P�c��KV+���!2��\�
�Tv�O��v`��VN��ٛS=���T��K`+�Uo~����7�jU��~ҩE6î���rF�}ʀ�'�qEgS	/#�v��E�0�Q�)�4�1�0��~e�����c< ������U����r�(Sad���A��<R@6^V]SuiB���Db�J�v����e���VP�.sJ�����a����pa���ZoOi�RkS��'��5Ea�
o���`/ܭA+:SfU���>�'_j�:1�mJ3���u4;w��k�ӆoNu;ٶM!����U����i�޹&�\��Zѩ5+���0{�֥���J#�?���)MSw]�6�pU^L��m��Ty�K/��B+�CZA��4�iO������#�&��a=ZE�2�q�*�����ړ�U2�؜6�,��|�j%������ƽ���^y���S��Fn�w�;�5�W�����e�.��}L/����W�����/��]6]؟|O�n�s_Nm�Y_�K(��q`́.xj\��]��ln�c�!c��<�M���>mǠs(�utn�Wֹ�;�K6�8�Ȇ*s�e8�����9�T���.��Z�W�2҆@d^�0 ��u�0dv��3�����+^��4(�q��<�֠wg�p��M��`Oּ�mf�/�~q�˃���˘�T����o����������CR���/���6_�w_ʏ���O��ϟ�~����PK   �sX��k��E  �E  /   images/022bbf54-c303-4c74-b4b0-cecd35afa1b1.png 6@ɿ�PNG

   IHDR   d   �   xu��   	pHYs  N  N���   tEXtSoftware www.inkscape.org��<  E@IDATx��x\�u&�N/���7��Da)��HI�$Z���e�%�ˮb����'y�'�M������v�8Jb'^'.�-[���(J")�I�$@�c�����|��p ���x�=�s�ν�|�}�9�v8�|%�N��؁pm-��(�ΝCa_�������4�Ʊ�"E�he%� JN��gl�k�ą��|��X��AF#�M&���/����)����o>��~2��CB���i"�w܁��C�O�Io5�O8��� \R�*r����p�����v�	4=�~ǒ�l3MM��>�l6�WU���sss�D�> k0��_�2�?Beeh(/���bQjll�S�<��P}��33�S]������m�����҂��wvtvv��ѣ}�[Q~�8�rr���t۶m�1CF}}=���&&�]q��!ozȄO9�_�٬h�?6n܈2%H����m�f2�6~��qL[�E�_��ŭ�78���0!E�m>������4��}�R*�K=6�iΝ=���dv����ON���`t�ҡUU"�w�1����#'IM:
���!�j�
��i���"���$�M�$�%���ۗ{�����'Ω)]eU�>L�pz9�y�4��D"���F�7^��+p��W4�b�B)���b:���J%�,����2�'�y�O�1�筧Yv�JS)84�%��S��� �X��S�ۺgJɀz�����p�"4�5�=�"�n���Wn�0�� 9%�c�M���4���W5������*a�ܔܓ<c.|��kQB/'5<+m�˅�O��N���jkCKk+L���^�!�C���nA&r1������~=���~Q_vN��GE��ϫ���P�n��W0��[Ք��]]�纪�T�ja�SN}SZ2�p6Z�zZ%�ד��Bd!���_����k_�����&�!"5}�w��������7uB�#GPH5+�!՗}a�gΠ�jtQ`���]D��k�~{�	�P3��^z5bCR�dn�Y)!����o_�*u��:i�.B�';��څ��%|x��]dd��O�iK�c]�!�.�a��Z��L%����HS"j|>\�};J����/߲���NFQ!i2i�3V�*Mfe�<��?L�h�狌�����1����^K���5O�!*��:���-H��y�5��Y-6x�N��+G�3�Ty+�6L|��l�L0i���ʎ4�6�gi�m�(
i'���
������x>�\Ty*3�٨沮���0[t@�s[�����W�>Q�C��0��(|9bϐn�����r� ���9a��5�7�N!���^���m�q�p��X�b��j����*�"���x�4���8i\|]��Qd�c��|y��͟Axa�^��$�IJ��N�bnaɴ.+&�#�I�-��_w�z��XM���Fجh��\��m{��L�'�r�12��z�h
F.�fF���yas5\�2�ӫ[e��|Y4W�S22���D҅������w�Ygh��FJH��E(�D4:kx>/��b��.,��H:m�]��ɉN-�vy0Oc���2*�ބ�[���G�Ӧ�̃r�G����܂gE��,l�ڼ�Z���@o�шC�c�Z�����ևR;�������.#)���]�
�eɚ�&��$6Ϡ�ʅHxv��x�T�f7m^�``�ΝƖ���\S�#�9��/uIaZ�5z3^/z?{�[����ù�]��lvgL�7Í ��Q�RGb������i�0k}��V����?�s��&颦���{"�bw2�-&~.�6�}��1�D,Gc���j
s	��&��6;��G៞ŝw���q�o+�~F���Z,<�0RP�����vh��Bo)ΈQ���	m1�c2�F��)�3�f��_t;R��}wG�_���3�ޥ�,7Ğzmi K(��;{�F�A�ϳ;���!	����D9R33 ]j�|X��-���IcW15�W7]���:�g�(.`� R��*����.���btv����8�;�(��Eȵ:dBy�:�S%��z3�"�'lhlZ�P(��~[�lĉ�Hj֜=F��EE�p{|��X@k�Eث�`.*R����HU��,L&P��K8c߀�M��;188@}��$tOs�ԔsA?2)+�:~�sp{�.3�kq(�g�����,u�����ux��6W���Xq�o}�2�4�r�2tz4j�M�-�~�5�2�8������O`��6�iÅaV��O�g?S_hrx1�����m�v�����{��4�i�"H�KKf�*�"����:ׯ��A������W�4l�$��]��8=ҋ�(-,C�Z�d�ʸ,�(����!���ވý	,0�3QZ�r��_&��B!=�*Q;a��	9Qå�������+I�le@e��0��#��kZ����Z�<Ȧ��e��(�zG>Cd�..'D�Q�S�#��#�a=�"Ex,��n�R�'��
�e�F`h��23�����>0%7��y�ٌ���k	
{����f���o��b���ލk��n���=hFƍY-�����TW��o�e�-��ɒ��%����:G�6]�[�~�Z+*ࠇe�~�^�Dq��5%4.&$���1ڌ�c:�T��9�xtA7��R~٢U�U?�B!=�>��<��1!�޺y�&��b��F{���˺/����XX�&���!�̫x��l��ԑ8�`s�y`�%��p���j����go%f8k���Ѻu�g#�ɱ�Z�)�̢�h��RN��"�n^���ڇ U3ccx�'����gW ��,�{�1lglFWeCdv�����M%�� 6F�=���1��@8m��Q�G�ըu�p8��G��)��y���pi��jr�a!GCܳ��T`rj�?�8
8��^�����(�l��������vS|�I�����:��A¨�BzCK1n�[$A␫"��>��.k	&&&��Z�C����*�*�����}��1l۽��1�]���X=^��X3<�VS���V�R�tv��ర�иaM�t���O��?���3��S]fך2�j6��w�\�K6!�MKVze�R�`&���H����� �����S��؜��T��a����={�־�����.4>���eed�*�Ed=�X@��P1B���엋��WXT�L_o���F�S0a�,�mi��{��������u�pӧ?OW�~�:�M���<\��=��$����O"I3��	�c�ԛ�ښNS�P� JOK�¾ibƭ�f�������_�o��ޱ�{�����$|�lHI�T���0��5��*�u ���_�6$D����?�3� �Ŋ�����8u
Z^��,!��/,x�h��)̻��j�d�QN��rF�S(-+�Y�������K�;�6����VP�Ӈ��������F����Z++a���=0��@gG��[Ύ�c|&H�J�Ee8���� �q/�]��9�k������L���?tp4��H���k_�̔��;�N��������!T;�(���w���M)I�����n�u7��R8Lbb`H�Z�+��%^����+�12��D�?���_P*L8+��|���;E��B�\
�VB�/�t"g"����G
K��r��VZ
c�t �ԎYb�(Ecq�Lh�kq��DX�C�L�,�G�iC�1"?ӫP���c���@�KyY�[d8h�w͏ f@�����f��	(lD3nۢ�����f�^��&)q��0�{%h�Dq⦨�4Y�����(
c6\�w�xT���	l�蒓&Sbt��b�c�[#3��E����t,\��oP���g!\z/��5�P�C)~��a&�pynk]��)Ӯ/�m؀�@2Z���ⳇA��hQ��h��7!�KOV�v�"�+���9^#��U�r�5�-�dU^^�.����	ÿ�5��x���0==�Æ�� ]L�z
�3p$f&�T��.�%�� ��W���������()50<c2�A�W�Ӓ̶��SmK���ŎYo�i3��yX�C(7{��SӸ0�,B,5��}�]0[97��b[%C1�VWG�F��T+��Ђcǎbnno�Ey ��m��ck�Cܶ�AA��A��_i7�4ҫ���� e6��]��ُ~��v�٘GF�ʄ ��#�>/�Jbp'�����I�C����<d@��)l,���*'3M/J����F�$�-��!D�s�|Z�U�<�8�)�K��r�r{�CC�3j��g�?�Fo_?:Ϟ�!\G�e`� �bXXH+w~>���\��#�i�7�?&8#W��3�t���-ڍtq12���$s�
ܖܻ��ϧ}>Ȫ�Fz,��
���8nܴ�@�AuMM>̓I�sNµ�l�c`hS�3�ÀpO\��2�B�.�c%_���BT��쇍�zyפ�H�CA��$+������3�RQ��E>.�s&#�S����遚�n����Re��G�m���_���tm�ˉ%3�f��g��27�!6 \���͛�d�/\�C@F8�lAICJ�=����TI۹s疁p����*n�Yl�Ԏ�pM��2���V��eZ���'>�؍7b��sϭ�A� M�5���ʠ����
���EY'9�Y ܰ
�=�5�d�r���s�Al�UA�����"�>$��Ӱ&�JZp�����Ј����d���2�=5�ɲ1#�gN\@׬�"��5��"��}�D��J����YPx�DR���$�J��%s�����.A��������ضAA�1:'�:���	�w�H�w1��w1+&��Q|���}d�NC�"� \qu5/·=
�޸dRFn3/v�go�r{]�'�KJP�t.{�0D����)����|Sn	F�v��[��ŧ��'Oҋ�S`u6�H
��<}_�s��w�8UA�]QM!F��ɫ�p=YW2�h�4I ����)K��MQG��t��3��?��w�S�1��_A���N��f.A���'�E���Y�ut�.c]��|�4�%�ny�����"������譢�6�Y����{T�a6c],�߲$�=?k�� �W�p�ٓX|W=�+�l�*Vuy)�Ʊ��5LLf��)$bs:�KQ5ӥcԛ0��v���Ipb��� t&�i�g��Q��/�C��l��az\�6��!E����J�+��n<�C \��9�-^�kO���ju�+�V�p���nW᾽��(/�������`�64cd6��[P�y�y-E�HF�29���,2�f��D0"Y<r�!RF�4�r�>�x+�Ԅ��F��nȲ�;���I<!�ԋM��u7ߌ	XlL.U�_Q�ʝ;a���0����h.��PX�S�
D�&��|xo��aN���L�R8���ˢ%!�T�=^���v쩪����@�nB[�m]�V�QWU���)��ֆ"�;/��E�`5��}M��G�U�P�f�����8�՞�4�:�-�կp��P˸��>�?���ϡ��@IC��ݻ|(�+wok^���r�[w^���u��@��3��F�r{�`aΒ�]wb=#׳g�T���~�R7:?���q:�k];�Uc4�{�6VxmFi�ґH��2
���c!����.�cw7�sg^�pSa`8Q�������e \.�����4��Ň��Nu6�n/U�>;�XZS�б��!\oQ1
�.�3*� 2$q�@���h�0��t8,d��67���B-�BY�2��2V*��-�+���Z���d82l_����z8���hݨ3��%�h��O�7�7��7�#�{��8�|׋>�p����ΉNGݪO&M	D�����u(E����/
�Ȕ����+e�I�J匵q6���aCMu��[yE9�O�.�p�dZ[[+lμ؍��z&����C�]]Іa�	c�zΏ��܈"GΏ�ctzAɌ	���#��?H��#w���D�n��~��o��y�E��"?Ĥ/��D*��F����|��M��&�##��W�'px��ю!Ը�(���L�y���,#z3v���E�$��'Pq�"��ku54�	Ő��/_f�s3s���a���AC�� �d!�1s4G)��)�b�NF�H�W��2�qῬ�5o؀-7�@ɗ_Ε.F�w�CW�K��b��$��Kq+&�ע�H�QY�G�ʆX,�,}
��d@�iz�Rɦ�ԍ/��c~L��&M[�C�a+
�s
��f�� \�J_�_x�*��+��w���p�-� r�b<��*��ȓO.:�	`�@�����"��]����Q����<�G3C3Z"��H���k*�89e�뼀�K5�pe>Iu�t?�;��yk�M�zN�6�X2�~{YꓩUoK�4$^�h�?�c̈Q��^���"�3߂��.�f�P@��a�.h+Pg�Rqxc̛��d�p�E)a�;���ő���p8���l*�ȅ[�4�H}�?	�ê�p���$��N��YXb�0QF���KW^�C�x���/��f�B���xQ.�.]�,�;SX�`��%S�#���NY�'sƩQ��u��E#u�Ӎ�D�#���Ae��%b��@t|ե�[��WU�[n�&�����&2h�L`[�C�Q���!�!ѦU�m���t��ѭ���QB�l�ַPt�z/�m�����E�L��N��	f�VU�Y���wl��.Q�440�ym��+���Ux׻�?�@_� ::�*׾­)�"�!܅�6U9�{N�d�ל|����ܚ���{/��mN���H �ZD��<�l�*��Ilh�!�B`α��Ƥ_ ܷn!v~�{�$t��ֲ���N;"zM Y�W�p�!�ǘ���s U��5Wb(�;G$HiF�~#7M��3୹����f��2JKJ��q�=�D޵�-��,�� ܎��t���p��Fsn(S�����!E	�#uIa�z*=׍W�Z��ǹsg��e�uzT�p=eh]�C�[6oDg�(��c�U�
۱��K����~����x������44_C�N�e�<�HX��\�`����6on�kݓH-�pӌmd%D ����G�`��0���q�vˡP�@�������*�HXes�`N���(�͆�N��܌��K[֒��Lep��������H�B�T߬�q�#�����4�F������:�t�(7i@��$ʥ�hmi�J_����'u׵o�*�VIb�%���P�1��#��0�v���p�
� �y��e!\��W�4�kVK#Z�Q��/�j�W&�.Aj�p̆��(�V#c�!�I�W�jx�� 
�nX6�ա��p3ٕ j"Ix��QP*+�ѡ|p��F�F}|lZ�CLYR�/�pm^x�k�
W�ܷH���kw���.yΙ�Y�����2�vH���U��
ᴼ*\N��A����)�%ڨEe���o̔*��]�C�(齸�cC�$���W�p���Ϡ�*M�GTPH�8r����n!�SeW�p-�b���<7��K*�;�]�2��8�a	��s9���LF*��f �l<�MSeU��b��q	���cH��S�z]մ-iږ������`a�!tq��-t�T \�C���r��-���u7[�;�/[	�b���핕F��?�
����A�,����܄��0~����s���G:6O#o���|��f��(]F4%�K��d��A�QU�U�N9 َ�����I}()e��4x"(�Kn	�9WÇ��!�C���zL�Sx���]eQ�B�4&�~;v;K0=3�������nɃp�ء �
�^��%�v_�p��H_�q��� ���`��$k]C�0�t�H
���G�*�$6��P�.�)��P��z�%��Ǳ��=�k_���5����>��,���/"��/���{��yz<K!��"W����ɵf�Z����R����Q�c$c,� ��M
­p������CC#(��`7!��

��}--m�t}η�PN)uH�X$b,�K`(�����.�����pa@��b�xN��Ԯ�E8E"��!�冨�	e���U#�� [4�={�\�y�
�H��,G�-�w���C���;������	�*�e(_�������ކ�n��u�w��3�j:��?�V�YA���'���td%c�����ON^��C/ر�Y{��˭}��T«:[����~Y�T��3A�"�!\�͊��V�=>t��{�<M�D�g���$$ɈT�4;1ٰ��qx�7#�D�h c3��
Vb��Ao��i������t$�R4�i&*��%�<Ϣa��$�ܬ�A��Oo4��Z�ڽux��ֹ�P�v�f�U9w�?� �]{n�����%1�;�Jztν{U�E��\�Jj������A���h9��8OB&~��������h�\���B��d,��rkӟ�bT��t^xA堩�K�vY��J��U9B�׿ߣ��&`��k����`*i�`"B�JZsXUg������i�������d�y��mm�S-.j5^��[gV�b)=3Y8Qَ(J$�T�B�d
��7��݉����YLI�D1'/ݑ���?���S���`����记X֕a�.u!R�`�$偱(	�����2.�*��'�27�����������h��T �s���M2�J/%OlI�!r�tZ���Jc��e2�ؤ�!��V_I�ԇks�E��Q��1�����s����Z�S��B���I!�*�~|����m��L�3{�kg�p��+NN��P+r�Bm���"��'�F��kp��>xV�5a� �p�Rr~�!�m��c�,��K�Wc(����_oۦgB�V��'>���|��)ԁQ�mſנ�f2v�Y�#��=���ߩ�m݊��7�]��k�$������?��K�dXz�$9�V�"�ٝ$l)~���?�������R���/����ʳb@�O(����$��gt��q-���M���"ē��iz��?c�t��+ˎl����Y��������UP2
�k[y��cqI��g�������*H����[�7��� m��0A���2��ݸC4���ѥ.`Օ۸��M���Ϣ�=z�y�1�<���Zl���Q���H?��=~��|��f�r�!
���|�[�<��C���|5�`8���V����
�G�_~��Ԫ
C�^\v+Z�{q����w�]I6M��ǫ$�4��^}���~qDI�l�˿��R����a6�Mf��q��%�.���w�˅�ӧ�����������?���#�V�6t������wb�d��H0�ۚj����S�Z���\@bټ$a���Ʒ_ׂC	�ސ��n��m�J�/�/�V��;��d�/!ڢ
&�=18�����P����I���^ym��ؾ�w�#�p���q�O�B����۱M��q��-j.,T�R���U����S����L4������Jej����S���_������2����`~avw��C�h:�U����I(����Mz�$���#�ƥQ�ؚ�>$2�,��e�0d���d��K_���ê�Vv�˚���� -z��u*o�������3�I!�oO���ľ�B\��AxfD-2��:qvrN��YcÖ��g��6��Ů>L�Tl�J�ⲡWzQ�}E�a�n���\�鲗�z��JA:��n��GK���j����|��L·.9����_bڭ��&�����#m�$�-�������7�cphϽ�Zl�;ݜaQ�XN������5>G}�7�f��S���V�@�	�#|����^���͡CHQ�;i�[�4T�W��/|����k�y��ّu���-��/ɐ��HfH�A-�,�*����ϫ}l�u�Q�Jb�oVoc�DS�%���4'0?;���1�~w�8h0��� P��pS)5��͞������b
!�~��G>��N_~u RW�Ts3*}���vAN���ߩS:��!6D2M�h�tM]�<��݃��TȮ�VK���SJ�|%��(��l�9lٲ�S3����ڇf2-R5ٺ��C�=�U��mB@c���,Yz�eЩ��ދMo{�֌I*m�O������,5������g��&���ϔ��hz����]��l�o{+��F��"�z���bcjN��ޑ	�����I���.$W1$q���������J"���p��Sa�a?���]]������+���*������s��!;�;�'�P���4;��	<~j��̍��Ϟ�c&���P�5�T&cd�����a7٠�pC-��u7c������`W3��p�$FɌ�/��t��$Iv�a������ՃYbNd`q�0�Bߙ���K��]NݞH�&G5�j�MC2��Z�fC�$����콞7�=Pd,��bc6��a�\_|IS���|��}��e.�"וT7`:�-f��wYþ�������?�.�2L��ZhWD���ú�M���խ�Z���`����w��`NI�`S`��V��n�7�+#��	���y�&�$�QJ��`�-c��!��K���RAEj�7���'V$~v�2;�c�ܱ��eN�!��%�H��$#�b7�{s��Eydxe����Cx�LT����QT;���y�F3^(��]��C���x]b'��%�f�ͤq�X��v�=���E�?�J]�L���a�45^]CS�g�^�-�y�Mle%����*��/F&���<���;�����Q�LIl-�E{])Ο�c���p�{/2�7�a-y�4��_���ڵ�~W��=.)���JO2����H�*�jĲri��N�~�x�_�U%M�'遼��_�\��Ku�g2S]��[��ꨫ���(WU�F�TJG�){j�}��zz�Plڼ�^���D?��z����zFq	���Srv�����\�
C��C�i�����ٜ����?C�А����l�U�\�zPF�5S^sm)�iR�u6���*H[�&D�mR�o�7����7��뉊k�x����F���|�t�L�n:�#h<�
~����ֈa�)N��Us��P�"�
cs��p���x���}'�5Șlr�i�A�j�SM��4��� [�Zok�a�
X��65����1и[��q�ޛ1>>��f!���f���r�C~��v�z�"��
�b-��k뛛Q�	��D��e���^T�iS~?���)���Jc��WK��/F%{�fY��l�~z@umд$�XP�w��^����D$]�d��#�ծÌim��<K9���-[P�,�=����-���?$�6Z�9�����+�
R ����d~l!{�ʊn"�7ʨ�O,w�\�?ٍ�Io>��ꄖ�b��$��"����Gˢ�2I��i4��Ȕ&��!�!%ϟ���;��dJ5�p���:�g���=>���w��\��]�Ť��k0�'�����+U/ �;�{�����u�3[�Jq=�&��et��S���4��Q5��[��&�U|5���S[|�g��+��b���̻�Le�TH�-#����H5/�*E���Q� �e���MS�!:=}5��
Gy��Pz7��v8�����PT�Í�U�H�u�ѻ@��At�͈RJ�K��B���B�97m��:笕!�}x���曑s��##���_��M�k1ꢖT@�o;�ZXo/nel�<������z�Uܓ����!�P,(+t��6z�ύ`׮k�{΀p�­J�U���X��{1�j4T�
D�!�8�Y�?8�ˀ�jC��w�-�W�N��$|�j��)����-��XU�(�T�!��?��]�
�}��C�B��+(*�bbt���U�/N	
w͚���'?���͘�a�i �˲��/%Ҿ5C5�կ�F��{�A��ʻ����3�d;՝KjJd�CRl�[���L��[v_Ȼ�U����4�.�����`x�� \����{i���nF���E���F�˺>�$��q#<J��%����x���}E�t�����8RU��K��1m��uu����6��Tk�$o��1��K&W�pKUa��-�Ts���ڀp�Ce���
h椶R�,2���U��W���i�]�3�{[��1�Dy��6��V�̈́�;�t����х8�E���r��ń�P��vo�����A�$C<���/���a����Go��l��o}�T!���X��D��8��N���ؚ�p���ޫ6t	\͆.��W��EWW��]_��Ɩ��sH���v=��^<2��H%��k[l�4�zyX9	�]�ͨQQ��Jj�{0��ӢO��9���Y?��!NJ�!0C2j���pk����VS��wiS�< ��8�J�/!̊�0x���?�]R��Y-}D���avv@�D�>/w�츾ύ�5!	���Sp:,jAVr�--J]	ξ�Ɛ_�7 �K.��.�5� \9��H�Ӵ�r{����a�6���;$��?]����ʥ�p��+�W���s�n�"�.2�$��@ʃ��iC>�ݍ���С�[b�S����x�*�U�X���O�bC���\VA�z��^���u߲�o<�ASx?��>|]��1nI̠6t���������n��ܓ�u<��eYģ���"��r�ϖH��Q��gR����|>��f�6,��9�����3�ҩ�T�Vx&UޛLƔd8�.�m�t� ���Q��"����Je�-�ܖL�	��7��W�Ģ��g�]�r�Ue�P-}u�n�9J
l�'3����k�r��\6�\��Y�����$�38�uv��75�C`���9��[�wd�%5��!\(7�j����a&���PgQ�j]�M�W�.mY�Φu.βE=I\^�m��L�.��΋��j��F=���}�5 F�~��bF��x���d\
OQ���7c4�Q݀��R��sQ���
����ϪU�;�s1µ�R�Z:��<���)ع�v���T\��YV��睡߾5'O�X��򶤘�>�o�~;̲D���Cc� ���=��Ї�:v�%��b��&���)����7�lw�_�/��I����i�d��$�I����Y����� ��}�n숄q����'.�pݦ �� �t�b� Ji��Y���a}�;`N�����{��8�!�&F�ƾnBn7�T�e�G%8�ά ��9����Ke.ZHs�����q~溞l��P(����������4���/���+�3��F����wZ�:�;�����#A��$j%}����vԊ�A�K�@��[��6ӠW5T ~�_�DXM:KTL�ÊkF.b���PI	���$��Xq�bB�~P
v�)5����*����^l4�%�)�~�ս��8_�*�*iće�^��+L������ةj��x��LI�:����ʖ��v�K7ꒋŃU�x�ߎ]����n!2l�/T[�֭_�#熑�C�+�I|jh�Ցrrl��lgUF�tq��T�
]�d����!�6�̋WĨ?C�~���.Yf񼿸�:HW�Ӣ'ڙ��K�����D��4��ǲ�?/=g��3��-�}��追[[�p���bll3
g ܹr���	+N�a�X�O٪�p������QV[�zUEXX���I����a_�[�<�`�K���XK���6T��'�#���c7�iD,�����D�Ш����jI�cc��V�3�Ji�U1$� I���bh>��yz@7I��Ԝ��I���K�j�`�JA^�ق�9�=�9s#�>G;Y/����Z�"�>{�}h�я�����J�3ajZ���@��ȘU�-���T\'�8�����i1��5�xm����z���B/i���Env8,6x�[� \y�\ ܴ�_��,��F�mO=�Kɩ=u*�-��y�hT�U��s�S�̲�#�LO�eF�c�uF�i�H�w���cݽz�\�I�]<v��]�z��05��`-�*$9rrQ�Bc/.Bbh�}�4Yu=/��p�X ��ZǗ�et�#C��V9���39?\6��3;)	�����-���Sz����i�%���@'��tI�}����K�i�Nà�üf�}%S�ʅ�<=U��.����T���q�9�a��������,����
�gF�i;�WZOw-�dt��$��*F�N���5�.7dU�w���?����/ �ק�[��T�NI8*��jV�S�ɧ���YT�ژك���n��Վ)2���?9�"���/��u$���{`�Ou�
c���u�ۯC�U�ql�L`a�wc	_����p�j��I��g�E����"�������}X�5�4���\�G��Ɣd����{��#8zb3�2�vШ3R��8���\Uږm�i��B}��p v���GQ�@��E8J(ES�hh,�~:�k�]i�:.����Վ�c���BM" ���ޞgG�F}f��Z��bԅ����II�HF�$ >&�A��-�PluuzgkuQ���A����:f�2{~{��;�C�"�]��$��Fc�m�x���>�I�J��7���㊠"UmdN	m�����Ɉ2���zT�ZY:�9N�q������~�JD��õ33Hю��grmbEe�7wR2&\>T��a�ȃpK+Q^R�s��c��M���Zs���Xi���L���m`����å��޾���0��e�4�E)�蝟���6�KOm�0���,�ƚ��?��A�t�{q�[���� �l��p;86etwh܏�z#�)�a���3�A����nd�_�wd��?E��ɕ�c�F,қ1�$0T�
=�6h����NU�S�c�Ff��F_N�PI�L�K�=�R@@�l-��(6�G1L��iiZ������1����L�#0E"jV��`&���5��s���&N�M@���	�����!o��̕�CW����w�Sm�JCv�1;���Ν�����/D���P��W�H�0��SC�ƒ���C�aY���[�U����:�$�T�f��IǠ��%u#WT������e[�'���X
U��c��!��z����jxC�V��c6�7�N�^b�B}�Z�����q!������޷˔5��u�7ߴ���KU.�'n<�^�[�x_�d)U���Z��uI��Q(#kSKJPh$\g����"=��2גc���^�������wi>��Pn���E�~F�>���9ؠ ���a��cx:��� �*���<�#i�-���Ys!�(�"d���GUVz��� ǝ�ߏ�H?�����t��Q�|�l찳���%�Y(�j�n�i�6;f74aCM1}���Y��{�oü�pc
��R2��������k7����xyĿ�pE���o#CL�&��&zA����vȑc李6��J�ٖ�ȓ�}���أ��C-ӋJ�n�^����&'��t��5y��?�q줎�p�cc�:�+��A�.-���Dc�#� �8��ܚ�!E��w鐚��-�
�XM�h��&Qs�[l��_���q��k�JLB����}�r��d��H��pF�U���{q~��қ5��׍��.sE[c�0ƛQ%�.k���T-K9�i��mm�g?������X��'ϜA3U_�U~��!&�`e$�������lmT�J��:����S�"�a`h@����8zn	Kњ��ͦ�є��ob$�$ݩ�PN^�ݴl�q�������&�]m`�$$&��@�������R�}7��Q��`µ��\�Q��@��L$�V=���PT����֭��I�9���K)8([���d,�v
���:�<�������]F�#SSH�tW���V��T��8��q�4Ҥ9�	��YɈ�k�ذ3�-�Ų�)j�J�V����r�Ύ7K�E���R1��s�\փA&W���6F�'+�P%me��� o<�lO��:����ki���E�.���y��������;��g.�͂(�uJZ��3��W��c����9s�+��a���3+�,_�ޞ�q:�I�f�b�ka���O|BՇ����v��XF�$�������2j�
�!����?�3�2'_zI5Q����}�p}�K���Ҹ,�=�+�����K�p\]�+�˒�'�~�s�}��)!caȲ;��r	mH�����)���!:�"����|]^Ն��;� ���*���?�a�
�ڱ+��q�mHlۆ��rK��
����P���~;�n7���_`�l�|u��?�3�)4���5�}vі|oD�E��#M��=���0�)��U��k*C�j�*�y?�e*��j�5� ����l"���J��[^��'+I��e��T������l���`�ȋ�e9'��i�z�Q��lw��P~�4���T7�+�Z0c�͊��f4���oqӱb�ty�@k+4J���m�k��|�?D�\��ʯ|E�s��A��.t�Ch<r� ���V	��c�ފ�_D3�G�Q�!!��4rI�JGSS�ԇ����"�l� Z�s��������CSruI�J�%3d-)Kl��-(P?�m������A��I�䩾a���}�$B[8m^cZ�k�2�d6z����R������TY-N�>�̖-�#el!}kkk1G��I-4J�8(�����ΐ����~�X_���E>�ȣ�bj�.�>�8�y�����p��=X�CfdB/&r�9]�_�rie�5Y�¥�F���l&��k�Q�X���6nT	����"���YU�
t!��OiJ�v�()QK�Ҁ9B�/�9F�
�x���ݻs�%{�<I;3q�M�~�}�$L�KYo{{��g������"��(�CT?sΞ�>��g�j#��j���	*��e]��Bj�gΨf��晌���W^A���m�����2I�C��ke���u#���[[�P��QD��=�]�*�sr�~N�l���ꯎ�WҚIc�v�X��_#el'��x��H���y����d��(�L-��0^^
2�*\���Q��֭8E^M{��zzz0.]�8�=��Xm�JCf��jV"nY�MRuHR��a��t!��O�;+}�����C��6I��f��C�i�);Ք��]����	�H�+5-�)C���ڣ�2�Q��,da㎎�o���uQ)�Uu�����(���Cao$�"��4^O?'opͤ2��J=�0�7ߌ�(��nD�kՆ$�%U���TK��s�N���ܾa�va�0H�䚞��B��C|�0��]$�W
��ƵO<�Yڤڝ i\I��!�9�{L1N1�Aö���F��>� =���.���.�y�<y�0C��;����p!|zj
��_���T�YH���^%"�=	�d���c9_$Nv�\$F>+GiKވ2���˦�|?��9a&�6�.�K=\N�Hh�l��"{�׿�yzb�%��1�-0����!�Y�dw�)����]�Rm.,J��*��2&��M��P�%ILa�d�H.U6Nr�^�B���i����0�i���QĠЕ������%��\�    IEND�B`�PK   ��X���  �  /   images/10ca8052-f8e9-4304-b468-4eebebade650.pngmYeT\˖�����C��-�	��H#A�F�� �`A4��	���h$�C�p߽oެ������ڵ��kW��Ώ�FC	�
WEYA���<B��K��h� �F�((�$�h^������P����8AG!B}������?��#�P����?��n�~�'(?�!�_~�߃d�o�[[_;0���3ʣn��<�����<��W��������k�a�Z]�1�d�je����wIo�G�l�b�vvrq���+B�����2�+�����yW�-�0P���Aj�VP�'�q&��������`0� �+Ԏ�_LL��O�W@��1������������ȿulݭ�W��� +WO) 😿�߅<������O[������������=v��gy� 'I�'K�/)qM����v�ڔ4�$������Guqy�-������$��w&������6�����C���T��3�}C��O~����� Tdu�3�a}��J~8���U���NQdy<�ݻ�'���f*�fRx��n"�ƚ�|0�f�&�[U��w�Cg>���VLĢ����J�5l�%��(�}�9�0"��Hs�������~���f,�mz�Շ���&/�f�qiq�^���!�C'iO��A���,���ĸ�T�s=J��7��2A��;�=M�6G��� �zEZ~�y�}���+�z%��7%�:a#,��1���i١�2�pY]R�ʊ R D3hf0&�׌��*~O���F�֑�1�e\�᭠��gJu���*���?#������� $ =�e��r�V<��B7�P�p��&�]T�T�z>��x�u�d(۠�(��G`���B�hY�ۚ�@�4�<]�4)V�3CR�w���~@YE�9�|��t���Ÿ/�k���!x�2����%eͮ:�o�P3�f�
y�?�E��ݼ��d2}�V�&&s-׶� V4̚xStX�#�9�*+)��@2�pb�1�z�`)%�a�����z>���"^﫪^W�7�¹�\�{������x4�1LyC�4Ja�X֠]���n�����Y����Ɋ�m�\t=
3�)+}��5z"v!�6��0��,�j^QjK�u�g�I�I�|~�ڈ�z����S��6l��Ȳ\�����Z��$5%�՞p��Ǔ��cl-�t *i�M\|�C���0�	����o�|ߋ��>7����aؖ΀D��Lxu�Ve����ux��8�'���~L�>62��n�Ɔ@0\-%�E����*"߬��]���z�ƌ�Ӆ�4��c���M�v�����A"5T�H4��/�"d�4�N�ի���B�@N==�]�	����Pِ_�����$�T�Zꥼt�f��i�9��O;�>*�f�wa a���z"���	���/�~�Wj�-�P9O{1���;�l��p/ARZ������r�����(��TQ+c��z�Z�)��x�˵}ufY�����teN�t�C&��͙)��ª:퍎����We�~�!�x�+]�ū��9d6�Sy~]��h��qH�{L��x��7��8m2���y�$�r}q/�C�bg�����ʬga��LZ6Tdu�||�Mآ�IR:�k��Dx.��V��vK5Z�J㧢}��K)Ggh�Bu�ݒ *o��>Z<UQ;�ބI/�^a�Ѻ��yXƫ򶮍�Ip��]q�y�&p�'�����7��aϲ�_�[��؇P�p)k~X��sȷ���������'��~��������}J���R_V>BGХ���-&��RI}f?�>�A�3y��S�t�|�;M��;:䙼�����\��I�����M�o7�_[9�8UT�#L�K(d�X�e��z�bX�m!����\�ra�C�����5�u��-h�^��]�ܵ���h�ރ%}�̙�p��;��[�|�y��+'.9ė`�^y�|c"��#\QjL�U��d�=��A%O�v!�Rn��9�0�aL�ˤT�PkY�
J|q���).�Gt����9����R���$L���\_�GGL	�M	`v`��J�D�g42�t���B�V��WML��S�R�
,�i�j�B��\�I!���D䑇Yj!xK����ݭZʛ�h�����kT$�}�ւ�{S��F��R`��q�HwVs�bH���������U\��Q-C�yp�I8�\�>�m.��Ќ��ے����#a}_4�I�bք�����0k�}GoZs���Ũd�O�
�[1w�8��xXY����{���iN�?����Rrɡ�M��v���ĕѩt�=j��u��f``)��Ϸx�(���'�hضJe�mg�;8s�o���؆�2�&`��UD4�K!�[��쁰�Sh��T��FP�؎��&>����k�c �Pph*�M�>�Nv���6�0`Ԧq�9�k�sfX�YP����I�{�2��Wb}��*�k�	M�(��P`֫�����?峗_�7��S0,�Ś!'J1y� ��bgF� �0��e�-��q�ސ�Q�ь��z�*�����	��퇕x�xÈ�H�bs�c�F��?_0l�G)Pp����K���ϐݯ�����)+�z�+��U���Q���gl�aX�� 
�-nC�f���T�4�Ő����Ć�m9���F��eW"�O�_aR��P��1E1 r>d&F�B���B5Ba��QW�D)����(UX�%(��y�sH�b��鰓�w�OG���?SN�)(���d�^'X�����F�����Nԡ�F�J�m�f�����s���t�Z�r��0&t��"��<�9�~(Sc}��܈c`�!OQ������_\��;ޅ|�	N@A'!�V~?p&��d[������ԇf�X�d�w�*mW����I��h;����c?�õ��U��J��2o,o�,v}�o�Qt��v����[J�`�$��)�ΏB��.�V9�9�n*wa�,}q��;�~���HH	��W(�yc�Q��/.5�c`L���$W����b��#V��]�>���}�)��,_�?tH��+*�+��Ԯ�w�dx�ƆA�H��_ 5��yxd�x��$�ѱ��E�y��q��`	�R�^6pvw�N��p��&�f|� �^Z}�����y�_�SS�u�	b�,�[9s���X����*0ХM�62�vi�OMPg���!�����v���'�Y����*��t~\&u�5MV��˫Y0��
3����Q��9��䞶�rA	W���~�M�k+�h�^B�=&J+r<I�9|�¥e''n���υ�,��F�#p�<'.�hԖ\��߯���d#Z*>ۡ".B��O�3�z��vjw	#�+Tt�f�����Is*�\�X�]{������ϟǥ�:#�?I��\����V�qW��z�͵}q�� lޙ������-:���/���~�XG�aՕ�5W?�0�:��� ��k&�mA#_����0Oy�`W�s�,�`�Q�S�P=&>�:�=x��N�}�S����]��*��L�X�$���{�h�Z����,mwIc�e�<�rj����^��G`jHU��%��
�\4��}A�cv	�*�+��Uf��O��\����1�ʓE���(�I��t�h��p��V� �] u����F�(�B�]���3�({I���_b�B�͝��ʳck��]�_-���
��5X�+KF�[�;:�L�߅hT�&E� }F�its��_���~���-���/����\�
/��I�O�<Ƨ~@]�_<�&�W�)��RFZEj��1E-�J��_�9�S;��K`���Q����I ����5�pr�g���n�*�H�W����=.��<Uwn�t|~ơ	�~kq'<xP��`zEYe��R[ˮ��3yK�&>��Q�Ұ	a\0�~׵<Nn�밬
�\�,��Cp�XG��*L��Y�0TF��ؙW���L��6��RC��kh�!M�E����y	��ݱg��MC���LD
'	��n�G�n����^�ͯ��8����A!�N���z{X������;1�d�uC�6 =^`T�-�[j: }b~��}��ܶ�yzW����o<j#�}뙞��CeK���5H9��u�J�}�U5��A�O�:ffYE�Ռ3��]���w'��8�~#Z;w�[&T�H�B�:�A~�Q]���aZl)~/ګ�+�`����8>7Ǯ>�3�I��ٚ��Y�@VNL�'�M�9��*�L
:�j5�м5��H����§���;� �F�싒���!?R�0�f,c�m��h�.�=�f�.p���u�Rnf<�Oݣ���`1��g��(99���9��;�jTf8��M���ɴ�-ɒ@Hle{�}y8/Ts��e���.�W��7���4Oi�B���n�1�-�O��\;�M�]���.�%�/R������8a;^Di��%b��ä�2d����-�@c�$�5�͠ E[����+��/Bt6=�B���c���1�h��G��nY?�%��E��=�iH�غ��mw�:��)�v�0�ވaCb���J#���E���@��ڍ� q[V�����s^�}p�F/)�	#c��pv�ͤ�Ly���{hz��9�dq;/�d'?l+�sJ춍�A�U�o墅�&?���5R�u~n�}.�Bd�;h�w�n�ܐBYc����XV, �����S����	ئ0�\�<��MP�^f!xz�e-��U�R;CE���;e��8��,�W�c�K����^���6Q���#p�P�QW9Ns��%�L7�%�^��IB'��^���zʔ�1�k�JW6�����@8�����������v��a�o�Q�c�:��d����#+�t c��J5׫�a�:z�[�-��tM�,	�B��'	1���ٮo�"w#+�P��⪂[�Fk��jX��"�3���=����n�߿�J�P�T܆ֵ,yԝ�&+|���¥��q���Ň�ou��;��/N9n'ە������U��r��)sX���p3��0{�a}��j� �\y�~��k���Q�����\ɰg�8U�'@!��~��/�G���C����^��\$Q����[�j��=��,l��;��ɫ�q�F��[��i$r?�AU�PRb��oxG��}왇��Δ��?	-�`lhq1�#G�A��Іq�K�H6 �L�e;h
o?�u���?ۧ�٪���q�j��TPC)�1�@U�Zh@Mǲ}��d^+a��x�3�g��n��m�qh	�4��b�NՉ3��q&(jh���羯b�3j���H�����{n����i�-��WC��w�ˇ�'?��x���$
�l{�,*GA�x-�����i_7��UE�T��t��7�� �[08'��2V�^���U>���s���!��c�'�2��Y�����k#���?����
�$v`�E�W</)d���>bGH}	s=��f��j�`��A9��g�a%pm�v|ad�3��ܯT �����-��%;I�G@�#f���L��.r�mHRg ����f�+r���;����4��+o�b�=gM6]ק;XdR���ֳ�E8�(�z��W���K����M���ǋ�[L�=k���9�Y���j����?�]����OII�-S�e�[ܦ9I�+��;���ۈ����	ZdJ����\�߇����xc�L#���X��3IlF��9���B�d�����L��zH�2�tL�:=��cg��W�T���؞m|���M�+f ��ǓT����;˼Aʅ��t�9=D\����V�<���������J���i�]��i�X"8�u���#2�����V	}y������MK�:���̠��ۍ���4f\$CHϦ2E��w,��H&w���[w�я��������gR]7��@ƃۘMم<���KjC�z7D�a��ey͚���Wm1v��+�T���0f�0�ੑ5��S<��Ӭc��ɲ�o}�v��wP�r]b��p�,<��1Y��ߜz��^����z���%!a�Ԥ����x�����Z���pO��P�f��D�\#]�ՙ�Ҽ?-�B�2.5uE'=:l�zt癊p���#W�)CK�s{ŊY�ˀ�%~�Ss���
c�����e����팭5ޖ�X�&e_�R2V�<��D(�`T8�5[m����B
��~�.V-l�H�ʞIx��k�K�Y�'M�@�?�����W��*��������Č|;�g��8���"Bdc`��X,��uj܅��wrd�h�ӹ�6�{��K�a����p�@8?/|���i(��G���&�O��y��Y1�~�㷉kKmU�
(�Þ�8}�Cl��)vu�d�(�jDj��q�sz�d�ih@J�ů�]��?0ڄ��5��#��p��R�{l6�4� b�L��JRSy7hU|VW�T�4
j%+ᾟ�JD�)dd>�h=�'���o��m��0��]����MRV�?�H5�F+c�
01���4�V��.5.//˽ta+#K�||M�11�B�gJF��w=D"հ�����6o>}Q��M)��憙�Ȋ�)*ɸ��?P���?g��՛���i0c�!��,E���x�$��3�0�i�կ�ค�d}�Q�Љ��C��\�`QKQ�`Y$f�a�����fWne�}��svZ���%���/���km�'�6K�ӳ��+:��L�^F=�k�9�*+=-�J\l�k��Y�ο�o��^���ޥ
|v*Lg�o	���ǧ�3�<��..��y�U��)$z�7+z�2�O���\�Í�5�5���*�Z�3Q�ԛXc�Hi���&Y��q�v��'%�:�bU�m=T?�X���,B�WQ�F ȡs��R[�s}W-)O���+��vy������a����PJFf��2E�B��OR�K����N7����UGjB�{u�	�H�\�*#);ì�������5�zz�{�hWK�&Zm�t������FO�*_Y��J����_o[˱-�G����8b�����.w�lW��r��`����]��s�1��)v�l�>_�ͮ��*pj�L/y5�_�����G�hG�n�8q����3h�XGy��T�>Q��X��ț�����(�"��Z���� �c�&��i ֕Iau}�M��{@����b�`B�����t&��h���U$w��V�8	V�l�k?9�U���(۠:r)�FjcP����v��O�W���j�a}�����{�uc
��d{�������']��xsGk����g��4ĉ�r����;'_�Z��B���>�x�N�2���ݦ�������������R��A�='�t�S9�I��=� �v��~����j�rQF�ֺj&��'	�����|֘�2�+�: *�t����J�xW�����s���_4L"�$� �����܆SOTS�٭�<KI���͘�}*���g:�:p�@µ�E��^�[�
&����~����k4(O)'�h�fT�X�=M�d������w��r��[�����E�ˀ )**�|�q�J�
�2�hW�ۑ%���:ڥ��p��@�垓��[�� �K~�%�����*y��v
MdY�����RX�zz��v�c)�d��h/����7W商B����PK   �sXUs?��B  0 /   images/1e112c27-401d-49ee-8ccd-a7b22cee0ece.png�]	8�i�?2є�LJ��]	I��F�!
�-�$Y��XS&�QيPd=�z�#�F��������~��4���f溾�.y�������w?��qR��ꕼ+	�j��G�	�k�:�l��㻟����p\�
�`�����+��!aqQ���n��m���^�#5���5
�X��z���5��o<��J,�t1���y�'m7v��ј�o��o�O)���vފ޴,"���Vbۄw�T���?���;���|s7�F]�������7}˅�㬺�̺)q����Ӎ
�<�ȓm�ޣa>^J5��ؑ���_���PX�4L�? ������@�i���ٹ�tΣ�,�?�)5}&h4Z���r���G(Seb�ӣ�g������П/���,�^)�s��i�S݆�0�v�Ź%��Y���NI)xϟ��ӈ��/�t�vxM�-N�*�e��888�D6��}���4�Aia����2�T�=��3�?���Euu5��5k���3�:x���t�P�X�k��p���JN�a!{"+�mr
�ƃõq�)�d���{�,�zs2f(���2���?M
_�4�:Ѯ;#j:,��{���/Ve���RRҥ+R������-�Ԟ�C��SY�9/zKKK�PUv��L=�(�`E���X��ׅ��!.� Z���ϕU#�(<��N��l�Slf����g�o�F7�>�j�v�0�0_݂6�p��ɺ����k��)�����쌈b�A����u8qK;`��'Y�������z�����E�{�1-�ڡŎ M���y�
[�验�����-����0�[�7�jse�:w��f��:3W�A�ޓ�%��];�)�hП_[�c���{�a����T��s�WW���8܂�=6n�"c�l�`u[a�%ɘ9��:Y�3�����1�6�i����pL�u�Պ�p*䔢o�B5��gϼ/���,J2O����s\�?	'�/3�KJI�Q�G�yë�~6���͞�HKK�\3�5���쪴�!!��1y�GC�Sbqqq����㬾T�����ҭ��u/5*x�����Q��/�z��G���Y�@��800Pc��;� Ӏ�jw&�]x.���5;� �-�z�,)k�G|�I���������*���w���#^��pم_��vZg\�f�@_�g�w�i�׉��ǈ�c���SK�����3� �{hq);�&�x�*�F=�uFD���9	����K0�\��Q5a��_߲%������cn|���}1A��P<�D�!R�n�>gA.���J�T�����::FC�	�	���R�s��3򿟒���q7?�`-n����2~���ʪg��Q����.���a��T`)���-����J���G}3*j��v3g_�ܖ�l�����'3�>�N����<�M=[%��0��vj�$o��lL���)��љ�A�m��;+%f潣�3�o�yO�����L}
/Ӏ��J6�ˬ)���u �JL���jΒ��	i��$�p�!g ��3��~ #f$�uйm���-f$_C�pW�f`ه+���uI�?�̉>"�=L�a��u� k�������YM�x���3�0�򫓞:L�vu�����>bL#P�zcIz�-R����Oψ,���7%:�e��y��WR�0omO0#l�h�v�E#x+s۞��l��X�u6b�<��)�.�U�d��^}t��ǘ��r~?ć��>�{�8�E-��U��F]����YJNn���/eL�9�0|�&Z:���n�w�9���[��t�jln�5*�(��֙�ǵ�5c4=��iJ4d�?A������R�6�x|��HQ�Ϛ�uJ'�:-q�m���'�YFtT�Gt��s;�-��|�?�I&+�ܿ-_� o�(!3�Z�[/]���a8�r^�O���蛈j�y�XQ���j(� ?���8��i�(��g��z���g��k�^�8��jA�tz~4�m��23����B�Sjqk��@�=Q�1#�p�!��o��w����5~���!����LF:j�1�	ߘ�<#�Ttt��s,_���� �P-4~8Z�ؔ����b���1'�����<*ϩ�M'�
}�Ɇ��EP�Z2 \{ؔ1���.@'������2g��g�B������GA:ӑA��\q]�$J|'T�ԓ��q��T�o�6�@9w�p�8���B_���)(Ȱz�����$��>=�jtI|�Q-��sn����x��2i�}Bx����=lchEI�DTv]�4H3�}o���@.�e�P��?1<���,k�5Z��5޿:��p"��bQ�q5q�}3e�C���/����/�����d�/��y�n9��%��A�4���{��M����x2(�l������Q7���b������	'2i�i}t��`$ŖS:���=�H�b���/55�r�#���Ā����M�i�6�$�V3�[#y,x�n:�GF|�۸�N�yzz�'�odr�bi�x@��ڙ<_G ��o|�v�[�����m�� ��Q�aknN��G��y�yW���A�����g����F�;��W���D��W[���|ƌ��@�MLL5��UYl`�bw��4	�&[Ɯn���/�������u��T�J����+��!r�_)3B�#����Oz���4�X��m�W�q�U�
�vxƈs�fxC3pl�{�[pR�2�UP{y�#�b�ȳ��0����'D2�w���\�T9��j6�_�]��&�|�朋�-��O���4���H]��:���ÌYY�����y�NDU͜�q�j��;U�7-���O>LI�X5b����!���(1]��X=������{q��79~���cx��ݫ���\m�8<��m���mJ�	Tve�@��
��O���w�N �*vLa�F���,��1����$o���j��,��O�8�_��!Z��#�!��&Y��b��ms��A4�LD�������b�#�����7x��5���X��^��/������Bo�Q�~ ���Z������Mh3�؞�@|Ճ�"M~/��c0����������½�g��*�_Ͱ�cf����pb ~)�)wv2����P�(����{+m5�!uC��>���b�w$t�M׏{���v2��m�h�,�ʅ�>�o�^2ҝi!�I6LSU��9��?��3����A&(~��
����{�@x64��N���P[HM"l~���X��]�ߠ�����l3�4S�3�����y��Hd�|�L>+�8�<)�`��1[����}|lz.J812j�0��P�2V���
�)�!������Ӟ��Ϧ�a�D_�_1�ȟ&.����	=W�n;���H�S��[;�V��A�U�G+�l�tj'�՞����n�_�;Ș�͋�]��u���e0�i�MM�/ �;����Lc#ڗ�=�Z��9�X�ob1"XG�����3j~�`�uj��7SR�������q��A��E����n/SR>KUP#݌W�����~"�洬n���kut��v�տi5�@����8�2~�����R�-o�)?�BiХP��}'Ӑ�9�IM��IQ�΄�}�m�����vFZ�Ӿ�S��6����6�Y������&ҍQ�P(>��J8m�[˪z[� hO��h��uߏ���h�!�B��������9��T0��G�,��x������k���p�� LU��s�������L6��?��w.}d�-�E�{��kq��\P\k��=]�����	mmm�����3�8ݱ�����4��� *�G)�g<���%q1��\*��T|�L(�tV�K�ֻ��P�)x��yo%�=V�� .C�Yg�����0;�@U��č7~�v�B�������C�rw9aا�0R�U�D	����K�]b�~]e����w�N���xm�b���2�{͒?�y�{u}��a���w������U�ǩ��C��i�z a����wo�d��þ�C��5�wm�$k6�Tn�ƽ���������;6aFQz&Z�b5�'O��ᨚg�ܠR�tυ`k3�qO}{�Hde���X�@��$� a/l[C���0Ж��ꈞp"��:y6�%�ma�+�9�Ώ���MלR�i�D���-Ï�Z(��4��I;W�8��	δ��
@J�ɿ8uj���}DE�\%���K~%�
�Yl������ԟ���5���4��#U�rL�y��0Đ6ϡ@W*��l�q�8�mV���\���ľ�3vx֏X���7��W�U�!r�;H`pj����B�)�! �b4�~���b���&������%'��,�O� �%����:�ĝOd���\�Ղqft!��f��y��&�\�^��Щ(�WgƇGi}e����/x�3 C�B3�'4N$���X�����������Ľ��&��:p,@�����R�L-�￫^|G�#�@	���N�
�T̣�х�C.|���|�ql~�-R\�D
��ot7LJM�+�nMϐn���C���	܌I�zs{ث��ӥ6�̐�Ԗ�1�\"-��D�m�5���Q8���f�����B��$���ن���j�84����ԍs�Vr��1bI�e)����xMm����&��W�N0�a%q��Hd�
g��-� o
%�~��'�����iM��zbQx���l���[�p։sVV=���/>C����IP��d��z0�f���8�����<全��M�7#��G��sE�q,�L�QN���4dlpʯ˵k�9��x&mQ�i�����^�C�ӌ5|��ꚛT��Z�=�;��Sv���3yj Q�)<�����9����^p��Z/Ns���^�5@ک݌�������9�%�}8�x�_@D*�/D3��-�I����l*��
ˎ��
���_��hE���M�dt��Xq1�
SB��[�S�&�ϬRv�|�3�����]���=O�u��me���g�6�8Ͽ 8��e���+2��sN!�9�o��{3(� �kI^C�	��)�*�r�����V���W�>c�R�р��:|��=8�����]�a+Ś׌Y�򕲫r4&��1�^B+^ ��������w&�z���L�cdҤ�|�ޑrO��G9��k�oj��y0�BS5�����o�N{�l� ڀ�����B�J�����,�'m棘_a��R��7��97��G��'Lԅ�:iB8z?"\�ÿ�Ӹ�X�C��y�֯x#D*�h����v8�!?�	��z���uL^���:m3�t����1���8��XoS�&�r��}*[�tmE������_�Hj8��:{N�_�y8�R�u��e�����
����^uoN��7�%�ψ����	'`���>
��y6�<�)5�-b�a,�o�rl�M}�;l��a5�UD��i�&����2:*k������̼�p��)$�ٳgY�1C�Nkq�DZLCH�l��8��l����^`����A��3XR�i"��@U:��B�;գ	�r~%�?Z����&d�-��>RQ�(m�%i� C�^N�ǂ��xA�n�3CQ��8�!K@J�����:FN(����&���*��;ܱHi<���bS�c����Nߓ�bcy��cZ
���y�k��� ��E��s�ۊ:���̴�Xɳ����/�\e3o�����Pf�v����.���Vkj�t*NHU�Z�$j~��nB�6�+��r.Ҫj�cku�O���Hb�3~�R�.�X�2�ȏL�?� '��Jr�a��ge���#6ŧ~��l��A�. �~�r�־u��L�t=�ւ����� �!�E�3=�V�����O�G�� ���$C�{��T��(i��;Mb��x�p1��M+&DbZ��O�ߘ3V�M�s��W�l���o'���*�L����铷Z��w�s����쎝�	0����%��$~)������ �ہgA����P:���ح��*�R��\t����q��1���<��P �l�����4q���Gɮ5��;�H��Rv���K�X�bzu}f 5�l8u�<UU�kF��s�|F4rq�f͚5^�� '���bN�Ί���4˚��)���S�@��s�̀uڡa!�=�&�xDw1���X���'����G��J�M8�7��L����p��8��Y��D��|fIj��/6&�2�)QO��l��&�<N֌+_XX��YH~?����<-��榦�)'Yr��G�)�Va1�lp"��(���N�p���Prrַ�IWcē*���ľV�%���ش<�dP4���}$���ͽ��u�I��1��x
N���w�&5�$�]�p�Ps����O�5�͉\=���O:�k�� ���S�����ƣ�N�J42+7�����jԽ��bdj���Q[��䶶��^���l��Gݞ�
���S��-,x�l�7ߺC3���c�VUiH2+�{��A5o{⻀�a#��ST4��yӢ�R��H3�D$je�({};�}k�a"Î;�3�P�uy^�Fiq��ƣB��T�0����%)�]II��;㈮k��bh�oi���Sؓ8��>�ۗ��*Ӄ6���͌�u�hج��37�(�>��9�s<&F�J�����c��b�k89}�2p"j�1{��=?��}��,��eg������?�!�c}������7ïSu�ʪ;;;�m��3�)g5��8!���e��h\�Йk��g��M�a� �+��Vj��߫d�i�$p�F?�n ���М�b��h����D�$�����`K=�%��2��!���9����P¤B޳��<={�}�A����`����`W]��98�uvP�g����bIa�&�S\P��:݂�X}N�}���&,��N�p-d�E�d�0'��pN�8������&(��~�J��4�8�I�Ȉ�m@ii铝�3��E�I2�Q'��u:һ��%qp�ōF�j ��v��8jq-�K��I�Qh���G��b�v3^H��9uІ�119I�:�,R�+�ly��|1&��^#�l[�0��Mg4���f��S�����]͋_�1�}E��ܲk/�6���<y/�S[`��+:o�I&��zH��#,�'s)��)��X�����oe���Y�'���j>4����(�>^�; #������F�4�p�wrL�@oO���s��������oM�b`�[�J��e/	;r>'i&�ݩ�����|��H/�+��F'��GhϜ���!���C+j�*��W�D���YG''�������r����h��Ei����)O*����k��EV6�V�Ei�[��*�>�G(�nÓc�����ܶ@��Cy0_��T�	����M"�3٠��^OA���}���3�T0^(�=IX��^�k�ͣ���vW��2 ��LO z��=���C����C2l?���|�~P=�>FMv����X(Id�o�F�{ץIu�jL3�������u��ƕ���fkQ<��F#� ��)�-���B-,���̘e�mI|��a�.��gϞ-�=�$�'���j�l�A؉k����8���sE�$
��|�J�O��,CQs{{1()�ui��:k�:;��D�p���\��
\5���\o�!����)�̆���v\hm��������9`�?�e p��*'k�t�F��^�%�-�"�I��*�%!���b+�)��g�/�a����X��y�,�����������I������Ċ���,c����;:L�;��>����l���6܀��>�ى����3}8���?P���lR��,��y�QIuΗ��k@~�fу@�N�ģM�y�ٕ�@��(!�t'?|�6l�����{Ow�@!Mǹ��(�.(Ř]�k��M�[~����;w<�b(:��3�p��q���Ȥe��G�#_�5:�G��I�ΗJ`E�JNaa,��^ZG�v��5������`������Wc^��sP��������۸K��^�� <�>��
j���:X��l������1�+17D��l�K�Х��bC�9!9�!q��^��M����~Ţ%�q�N���:��.y��~7CX��MsH�.(1͌�;�}�����l�a��8c�����AFz�,Iw4�A�f�����Q�1����ٟ�\�w<N�k���^���!h\��F����"�������V��ڜj�	�k()����B�I�`��,�_��c�;�ev>o%��05����2�ste�n�YU����h7
�a��'[���M�d�G��t�<fn��w�ͷ����M�<���;��Q�sB��Yc��SC�<�Ucip�,s�b��[ۯ�X��b���r�S��@���r���::���ۖ��۲��M�s��_�ѡ�����7��ޭaw���6��P4��t�'UՄa��F�����MD����Jk��>M�:rc%A��dUS *��e$f �X��69f���$���@٦���ZGcn�:����FP��qXX	d�|��M���&͡��RL�{�x�;�ܖ��C3�{�t��S�m�ǹo����
��]��w>/?�pǨ�ퟟQ#g���w�c�W�_0�r���#1�'��pD��%�����������õ+F;�f?,̡�.�Z��f&f6%JⰪ[@��ܸ��7��۬c"*-�e4�����`�X��'��[�-�H��e֒��:Y&:gfdAs)��;XvY)�sTS..���J�����z��qFn�b��2�rZ�Nb,��ŵ�/��������W�(z\e�-BCC���>�c�A�\!�����=�L���k�OW��Z4A99��Q�Q�_"�p:l��!��b����#EX����A[a[����w%������$8W ��_jIBVYZZ&b���_�G��u_���1��'_`�"�{o��>;#�ܪ� �ȞV�tt�\�B㞪 !���9��Y����fAs��oV�ålhdT�-?x��{�$�b#���qq�@���+��C�p\/qY�Qbm���:zz�97�:��	��m@kU`
V�ݚ�8m������謗cDi��#<��W�X\��,�m�R�`n1����K[��y���T�T`�_��av_T��b�1-.-+l���A-=��+��U؎ ]���|�wwp�
��X�4�aYgD�_�+޻��R���g��Ě�qa��7j���<~>ôC����qgCc�rXt�ݮ�y���Oc�C\_��'��#��iqu|1c>mw��.�`*�v���������L���pUR���E�^+}d�w``�X��8�M� 
Y3�R�wmS��|T��15��h
�/������;�2"�R���5��#dꓞ�a.��8�T/��uDY4tN�
T�A�;�-3��sa�Q�L"D�
�r#��ZF�K!�S2b)����/F*]�8�����K\��5Fv]���M�y�f*�(0��9//(d�1��C���8)r����;��U`q�����C-A�����`>ٮ���h����=����1y����e�BRQ��@��`��a����$��|�i�J�z|�B홯vݏ�$��5Hs��~s��9#� ��bE�W��իW��	�oq�`o�{9f�icc*�1R�H@��%y���r8���F-99��𼃜��Gz{�u?�z5�J��abB�szkhW���6��]��v7��A�{��E}cq���K�/S+L�w��֌AY.a�1�eǎ&�
ϟ��;x�M8��S^C���j�[A�����4��S���5��ں.O�LUO�l캐��յ���K?�,1�:s�b�-VD�/�'��-:��
,���+�WS�M���l����C%�{D�,�wJbeM%��b�.P�5�[�e��^PT�����)�٭�E���mf"�aH[�����.t(٠����tk�U��%��V+��&.k�mn|`���<����8�$R��׫��8�󞗱7�B��}�˅b�4��"LO�}��h�Y�%�+�P�2��[+�Ǐw��������Pb��ll�_y9?����� �º:�1
�����]�3�^y�X�����'�R� ,���E3M���&;MA����:+� H8{�:p�'�K ����c{�Y��Te���#Ϲ_�
" v``|a�N��a��''Y�L���̀�P8�����<��=o�/S#�+�	���P\WyhJ��3S�5�%�Zض�3ֈ� h[윘� �¼<j�*B�i�Ue4�a*�w��o�����v����ra���lrF�;K���LM��@7�=�c���Zl����V�q�^j�8g����	�r��1@�BaI*
Թ��I����uuu��QU���p�Dޖ����H���sz���K����ع�]�_]����V[<��ׯ_��R<���0�t�ʺ�^I��w�<W�̇��?ڡ�|W�[a�wao�� �܆0�`�Z��tl[�D(��[_Z.[nn��΀Q]��\�p��>`�:�+�wS�.�P
=<=gk]�
8F����L�b ���͟E*����^��
���������i�B��T����zU�Fqf�X��0:*�=A�SF�v[��$oIƷ�*��K��(��PpN�Y��ICJb��M6���=ĂR�)+H�e�9k�58ɴ�2ۈ����j���� ��QI���]9Ȏ=�"��!	s��P���i��`І(oj��rtw�ihh �.�P��Y,���Yؔ��n`����3���`��v}㲟�@�X�	癠4!���g~<A�fqs◁����L��p�
��9,���Hn���6;�I�:��^�#W��#��3��q���w�" ��L.�FX'#��h�*(̫����L�ѧ�s�N��Ȯ�DsL\�Jy潕�{,��]���S�uSǥ�p��*���rj�?�t��k���'Q�Bk�9p`�F�wG����]�[���f4@M;��
�+XC�C��V�9ѯ�o��*W�����H��Im�tu��ҹ0;�y�R�4r�ŵ�S�Y����/|���Ge��	ʱ�n�$ܬ�7�7�l�9�Y wz^L��9hqZ�z�鹧-�ԅ4�Լ���6熾��5WB��W��ѡ'��.f����3�W Zʿ���� ���&��jDz�BB/��AC0��%8_�x���?�'����Z�f�J�M5���+:lռ�F���C�kF�$�A�=��3ǎ+�:��sV4Y��)�j9��/�ޮ��O���S�%�P�Wb�}`�ۚ�� �{Z��Z��,:�cN�e@���Pb�<N�z�W�U�_6��d�at�27P�L+E*�)�H����Áo΂�q?������4E��4����׶7}�j֓r�+�[���2���1�7�$u��Z��� "4|3�龜�XĹ����Z"��b�ÄY(6t�\;;������*_��>yd��/N�
��@�],+����p=7����XO�-1�
~��񐪜B�A����\kg��5d�����l,�����暱6�L{ H��m|Th��W��W�GSlB��"?��/U������x�
i�sn$P�bz�tv�ɰ
ٖϩ������]Z^QQ�������3�A�������"r��H�ߪ�
blҘ ��^o������pЃ�ng��Lq�[������i��Zĺ��L�9iT��5Xe�Q11sR�nNk~!�c�-��D0/kWХ���a�p���i����$�LT:��Yy�ԱYp����Z|�;M����a�`�ߵĘ�+���!�?�SKML*�d��w�W��ۙ d�1bR�[�*Z�pv�@_�8�5��A��3�� ��B!%�ƱP��|��-#�8��޺Q�)�~X�,㌄A6�K��k��䅅�)���ϥ�Kԏ�)��K}�g�N�%Z�����=I3�gI��rJFU����,������h�D�_���P���=j����\�~�W���V�ʍBõ	��DWP�^{5M��>�?��r��;q�%p:_�zر<ϱ�(���693}S��`�,:��lFQNA;h�bH��P�疶��t,u��}�� i.���@y�_N�w[{��]5�
}���Cv�x��ͮ�A&���� �e���


.��v�W��ر^����2�r�՞�æ��Y�C��5���B�BhC[x]�;�z���fLll�)���Sj8W&w]��*�t,�Cg�^�̫�		u�r{�}�l��Vc!��o�����/J/�����T����z�wF�b�9� qW<�n�*>�nyj��w�� DEE]\�Ueg�@G:�d�E7��8�t���(�_�J�e�]-��@zy��L���6��b�Ëqbwv�o�e�Rd��ۊ��?�:q�9W���e��o�&B������r�pX�S��Zn<�E�(�_����U�J�(�G�^�Ϻ�X�O"��a(��=i��;2��r�V�3���}�`���I Eފ�〞[�l���2v�yi�}��Rlk줢ʈ��H�x�'N9��zu֭�������gt��0���x^�����7��~b4�.R�&����I$RGLM�Х
i<���Z��UUU�+L�D����$Z}gw �sR�_�;�ƒ��?��mj�s����d!d�Q�QU� R��;�������Se����֨�#����m��� Yi� /�'���tژ|(;���_�Z[_@��\�;X5�S0dJ [��Q��ܘ���3�m	� ��\D?2�+g+/Hq�N�+ƹJo�ؕ��B�a9�L2�A9�.�놲��e�z�)�j7�"�K�D9�̓�>��V����k�+��b(�h݋Vx[)O KN|��C�_���ŃH�ϓTk�����_����@�j�E�#G�|�@4Y#�`>
��'���h�R��^V��L��������Uϥy�	2�5�wOvaE�*����+;v���Ӣ�î��n6�u�_.���X(�~H��䅙�c�j�--B$��`���1�~��]G��!�I ��&��W�����"߱<�e<n@�m?o�Tk�b��I�G���5��w�%l����?}�	�BjzQV���c3�n\fQ�tw�� m�Cn/�[/�*7���T0�*m��Cwԩ�h��$+�2d,�5dq;�C|Վ_�Q����,KE!�¶�D���E�c<��Fv����҇��t�i���j� ���~���#�L��mː�P��gD��x�lb�/�f�(�R�	���F\���Wa|��ּW��p�x�Pmg�ԉ�	�p��69:K�V��W樻?����-#�"�������.��2�l^`�咽*�Ȅv��e�B�-F�^���-E��7b����h�x���Gvm��(z���c����������������Q���~ﭶ�C>�)��ν)#����{�cN�iֈo��u�������4��<!�xg�V�
��ʿ���7�T_������_~澙z�W�M,���T>1e�v��ISO��q�Ě٭#ioԝ3Rj�,
J�v��伟i��I�/x�UN����������&������ѐ���$w. ��D����ጆBI޶��7j�Z���cd�hÆ��WS3�����\�"Hd`��F���;�.�^��E�{y�E�v�4݄Z��C8rV�M~��Ѯ��j���w�d*�3Jz�fG� zvL�0G�����\���f���V�۰_ɦQ�`*���z�~�V�8~7~�p'%8rѓ�1�u��w��J�����դ�Cef��N;��	���jڮ��-<�2�v�
M7��:J65H�@�k��m#�LB��tuY�J�|Ѷ[������d�!z�XP���j�2N�Nr��]\\��ͷ�*�{��A���SSS]'=���8W��E�y���v��U>�{4�NH���1;wțw��2�;�^�~-w,�ֳ���۵E6$@���0���\�pP�}Ϟ=������G^��/f���uꋷ�G@�r�����	��&b��Ŷ#W�0���m��]�ϹU�2��tn<�iJ�M̚C���D�h������8�F9��UQS�O����e�D���Aa�����>nli	����VM7HC�[@�%���~�f'��&�#�\��oJ����g�S%m��+�7@�_�  Wם14�؄���������/Ԍ�.��\ߞ��	A|b��3���=F���KEi�l`}ɍ���hy��3�-�8�����(b�U�`x���P�����h�q����(;;Y��]95�>��\�M7_;�K`�ޮۄ;ס^��I�����u&H7u}���sh��Mp�f������H%�����M�D�b�CN��ھ����h${|K�R]	�A��%�_���h))]Q���?�'��G�tW�^hlk�%B�Z�֣��	�;ؕ���=�΢ƭ���&������̙?��DmaB҃�K���Y+RS��|~j?��S�1��VN������3�O���c��2�*d>�vU�t���m�sn�j�@��-�z��I���-����9�������Wv��%�c�'�&��<���&�`��UP�HV�Cd�"�s� X��Vq5��@^X��ڝ�ON�R&5���������791������-���S�mꥠD��37]O�8������;^��������ڔ�I��j�l��$�y��aq99�����J;��M����������������ur��"�Oߨ��_v'�Fcss@���j���|�)��魮^e��E�>XKz��ڊ�GЊt�1_�Ϊ^��n�$�ir��k�PB���?S�hۨ���.9�8ϡ���'��<:clr��ZB]&�,��Ƿ�7xs�[�}����6R�����=M�9����q�}���My߮ ��i&�끻6�L��$ؗ�f'j�845�����$�~�knj���J�4f}4"׈D0�LKO�Z�/����֒����������Aj��� H �0���'b_<ȳ����6�^y0�iˀu�����S�'��b��KP�*F��="2�o�orv�vq���jBw���7��"ԉ�!Y�A\��Z{�u�)n�T�=K5���OA�8�ή����2�����?��J*++[�2���j�)
�A��dqk�v��@�yp��^58h����Uo�>�i�S)��� �����/z*/��}��szţ���W�!�§B��Ed�%�l:�>��_^��ٛR8X��{q�G	��v(a�$�:�`��w�p��ff�������2A��ܦIS���ݦ�X�{b\�s��>���Ǽ�=���+���B̭S��fˈfG��TPg�m���,I�У$7*#Ŏ�7�ʍ��{������|�Ւ�3���H�7v������ع�Q��\E �α�?_x�s����.I>4%�g5q�ՑE�22�<���&MT	C���,ι�ڻ�J��w-�6S�h%E�I����8�\�E;�o¾L[��\[~C��B�QGV��w��g�ȃ�o�72"6�y9� l�I���O��5�Y� ��fIf
�ފ|�'���7�cbb�b݌�x�Te�^�Ϧ�l~� ���R/K�����S�U���G�k��Ďx�W�e��l��`����m�e���t�;�i�K�fE�k;�*qN �$��GX��<=夤��aMb���U�~Ϊ�my���>
��}Hd�J��|�+��-�hހ�C
ѷ�tms�3�ȁL�����$��W?R%(22R��5iWp���K��^7%WP27�qɸ�A4�ť��T����>��H�#B�P^����9Gǽ�oN��	z�g���G���?(�$k��^h��<b��G_n���d���ׯ��WQ��FXF}�|1=�Kʗĺ_�ۖl�	��S�����Xc��S�g����iQz!{zK��{=�������n�E�|o/�@v/����t��D�_Sf~>OE� �j�(O���&��R��m$�^�)���c�QOH�B�vP�����d�J�l�֑~��4D��\g���ߵ�����{��!(C��g7��J�M�V���wz�r��/��`����kމ�f�{�d~��@�]�l�V�Ag����}i��'Lfޚ����.arc��>����|v+F�%y������/~1"""�ɖ��Gu���@��(��j���Œ�f�y�D)�o,�V�e@��)�d>{����@n1��}׾�'w�������5��-�A5ww?�VC�zpppcSӍ�G�/ �(e5\���bY���3"�#�Jl�7y���3���8�F�F�;��k���a
�*-����0�*�z��rU)�z%�O�n�^�N�M�Aл��L{]==�`Ec�	w��hD����z��z�v�� �ju�)�u��8�ç�H���O��hzσl�~� H<����|�5���~���q5��] '�b�XWhs�cIj�?����Rύ��+�X���OTT�o�@�5���׾*?�iM�;_>`�CO���?>�<��Rȹ]��.�������Dv�r�9+�[bP����t�����[*��f�'U���&�sa�����禊NL��(�:t�E�p[U�/o����q4�����q�pt�6l�`v�Ҟ;��?�,>�7��%�jzo)h��9	��"�ڣ�N�7��{/���"�V�6�@� Ā㧿��Z��HS���R��;Q�*���V~^��Կ�г,Iث���� c�jս�$/�Fi�]9`U9�L^����3,N����eiY 7bx�{�V8T,wgu��ę'PQ��x��$y�+���re(����I{�$Wrfơ����5��	0���%�J�~7=֓ �=Y|�`�Y�7��;}3�]tC �9�"����#CQ�_�ז��eZ�v�"Oc��d��E�8��l�! �Ʈx��Tʰ�I؎<���� �s�+�M2����?�c���(r���)�L�Ǝ�yo�
������9�E;�zo�&��:����$�nS�^C�s����^ч�����\"O��d�qt�.�0E�fEb�O��+�q��� Nq#(��GU�ɝGA;�%�L`��$��r���̧k��%���J� ��r���<T��
u�A �yZz#G|��yt��e ƹ�+Ȗ�z�A��}�3��,�M���b���⑁�#�PY��V�߾}�T��#�q�dU�H���X�㷦�O	�����O
>�iʒ�\����c�*���N���!��e�����;�(�&�|u�\䯁�EM��s�=��W��S�j��2�=Y�7��X�}��bY�]º�2UR�_O���C�Sܴ �j8�K��\�B �-���W�5�;�YV%=��|�~1]�s���Bğ/��$��R���d�P���7_?��᝗_z2��q[od�����j┆���i��I�l�{s}GQ!�h��ٞ;�K��H�D����bB>�qE��D��4���섹�H5�������垨����]k/�r�:�0�L��Q�v����Θ�&�j�~I�I0e?����q��Q<���@3�74�e*%?7\������\ٳ���6f���:V=��v��k"f�.+	I�7�(/W1,&��%E<&��{��S�F&":���5� �P#�������7�? �Ӣ��ˇ�,s4�ٵ��YKEm.��K�e

"���"TL��=US%#����O�3�[�)
>�Oxw�t��s�?�9V��E�>�V�	ɽ�mB�[g Y8�� +���u �� h����߂�#�	!��.��W��-i���j�|X"Z���mR��]x!�ê^����C����ޓ{�\�?��o�sc֙�gW�U�,d����W�ߟ�ۡ�6˞~z�6�i XQ3���j����'k$��T:Y,�ۗ�b� �n���q$+#�+U���q>�b���
���i;#-���-��AP�_j?H\�j��6QY �u2s'om]�9~c���y'	 h_��䖡��2�� 	��Εt�cd������sۿrS�;��@�����%�f�ZwN]�x1��t8���s������"�b����$���%X�GT�< ]
_J���V��[[U�����5��M&���@{��>'���"������g�.ZK��%j�m\��Hd�]���6?{��*�{����g���w�EH���@ֳg.W�v9��:y�w�FLX�nj����
�O��F�[Yd��{�uZ�&"�u�;;z ��<0q�ͯ�3l�c�3I�7Ͳ6VVVj=>�qquEL��-Jm�F��@辅��	�'X���Glќ�A���X��^-��m�#b�A��nD��Aϩ��JMM�V���*��ͭ�P���}M`Jh/�%�BX�xBFL˟�/h}b������A�=?B]�)5��\yl�E�����չ��18<�Nj= �VU����ŋ�N^�"�H����ʅRer���{8��t�|F�U�O�<�D��V��99;ru��1�M9��A�#� �8�����c����?�w��m�?9K���UN�v��Ҽ�HW S��/�(QF���}��� ���{K3��v�F�Y3{{�X���X�^�`'���5��UO�T߻Pl�U,}�����*S%d_��ےÿ�h�c��!���yCųܢ�Se�;�G"���fB��2��찖|m6�1?�
P�%�����q~֢�.�0������@���+q�yej��UT���/���%��&�-���24�'/z+=����
"��͞C� RR�����e�JF�����	�ӅmƂ�r����Zw���Uf5�d����Jde�k�w�MN�!>B�g�9-zȦ����I8�Y��D�����s�P�ɹ7�E�E����h��b`������nM����ɉGt���q�Z��{��DV�P'�{0k�p)�����M�]����L!6�C�vv���G��`�����oJ��FOG�tq
^o�5HCv�|�?������{�dC�zmj�~zqc�4��E)��0���("0�%B,m��J0tG�������-�zkQѸ��bQAX�`�	'�������m�=�1g?O�	���#�f�k�.��ov���F!���k�''"�zH5�+��^I �zg�;�;9�9���Y�wa�WA��Jq�նEzc<�,�F.g�C�[Xt��g}M��]7t���Җ�Lo2ɳ��Z��͖���YCdCs�)�6�Q!���۷�"bb��\�;��@uB��\�٦Y�޷au����Ad�P���*=E��������CV��D~=A�w�B���E�)32_E.�5�};F�X�ȥ�T-����r�b�k,�6�fm��A6�]�O]�{Y͊����V��ў��*:ѱ!B R�_���N�g�!(��ŠPa���4�G���ꖦ�tLW�ƺ�t�9�'p&`<#å�>C5u�hS6-��w�F���K��>'+�f�B��\E?qhk�U!�O���+��z{�����E�pK�"E�q+	�(�ʾe_��%�(�=�}7dO�}c߷�������~�?�y���s������y�s�]\95l֯Fj���W�������F�]%��XfsW�?�ӂ�Qʊ��0��LM�52��p�^w«�W��i�<[�rD1N�����7��7��'��c�Yhi9��Y��А���ޮ2F�v��LĒݫ��QKu\=������/�.�_ׂ��R�N�Ȓ���p��N��'
 ��=qt�Z��cp'|ff��Tw��bbO&4�q�1Ր�و�����{Sl���Q�S��Le�'��AlwQ)�$�oje!�4 Ԓ3�q�`������-�h��H�m!��� >��?��Z2���=~�'E*1�Fh��/E��Sq?�9�')�H��v��j¬1��^b��>y � ����%IK��˞�Z��U����vv��+��Xr�������Y	"τ7D�B%B��Դ��9�1+[�R3;Lk6��\�����*�L{�E�$,��� �����E�	�2(V�cb��&Pp���b�����r,��}�Ao�k�\Ib��8a��p��s��.��JΠ�?�{P��SR��ر���,s5c��OHA�Z<��LM>�Y�z?�E}�.=|,����Q<Yg3�8i7�l+鄍�<�����Z�p5%�#������8�2H�]��mqk׶��������+߭�Jf�rDN��,���iY�7Q�9�;����0��o<a̒%�C�G��gT��4���m�m��`x����}6X��	`.�� �{�b"�#"Δp#����j"�9��� rB����[ݴ�-�+�-�c<z,�{_r�9�M.ȡ�x�`I��a6�fYQTQ��c���e��ڃ��E���%2'�Pk�䴾��ꭄ���a%4zB��9J�C��uq�`4y�i�>�6�$�@)�!x�Jw�3�p_�Z?|2���_��ҹ](��p�c�@����z�"��G�7�0�-B�9�#nnn����V�&��gt׋x���u�s���zB����՜�-�4w[��b7ۓ��.�OmW�YD�ϙ���6�q.�w\9D�*�'�� ē�ج
N�nO����$C�n�,n�zM"� 媪���Du�gí�� *��$q��$��Q���7�4��^u�i�ˀd������i�ܴc!�Cm���=�F�����j��}�M�+�ʹ3\w*�<�������s������������.�0��R�nW����u�&�V��Z��N�J���pG����v14��ƒo�g��$J.��"�ep����k��������\��Y��ey�&$OBS2�p,3Z/��.N����Y�N���nf�ǵ�?���^�0D�l�N2�Ә�c��ٿ��A�1[�X��0�E3�s�h�>��\56��t*��]��������X4i8J�6%9|�����u�������W�u�3>���5���X����m^��p[����R!�3� L���y�1k�_~��x!�n�vK^ƹە��,��{L�� n���_'�=�d���/n�f���[���	̬����m�M�HZ��w�a���,��I��~����ި�%��� D���G&&&Z��U`_7���ܮ�o/,xyo�R�D�Պ��u[�$k �,A��k���&�h�]澡�����t(YM����k�>+��׿��vt�J�G-��(���o�r�,.f�^x
jf�8D2)�h�_.A�۶MA��z��Zb�e�B���z�����r���I��
_�W�)��ڮ��̵p����"&7E��/��$t���`=��lA�2ޞ�:\�5��Ur�M�<�!� �E�G�q���ɂ�M]"梩}��p����D�������ξ��rF(QA�o;�d�9Ӝ�Zq�ŷL&�M�k9�mm��ӥ�~�mNz�> kjR���o瞸���]�Vµe�C�ת*��K����y<`!�%I�p Ze��g��w(F��;�!u7L'r3<,K�B3^U�����
��Ř?�:�b�͛7x|��e�W�)�z@�v_��ͣ����,,,*J�O�����H$q��p�A&�<�͔���Rna�[\�q_MՓ�':t�t�^D�t<P�^Y�'��HsO����h��Eѕ��Oq���3��vB8ҕ��ᦴ�M�S_� �+H��:������@�6uޔ�����$i�3�Xi��eE"�%��x*)Rs}�ge��+6M/O�4���C{��6;	^����[��c\/�h�5�|A��߿��Ǘ�.��ћ�#Mz.c��X�ŀ�,a��r����Ȱ?`zz:e��%�WTT�X[�{U�<�"Q�������,^Z�O	����Ɖ���	��6v*��a����F�k#���]U*��F��-G/T=��t��&�}�.���
��������ɧv束}�6B�L�]#�ˮe�x�������zg $���e�lmm%$&�A�����K툯S~`�07;{	;�p��'��*ۋ�̀�<�������8�/`b�6,�O%�el�fT/���O.��I[AL������v�3,����0��%����Q����� ���{�#o�zzz�1�1��@v1֢$X����yy���S�j!����Ѕ۽%q뷩��y6�K�~�y�·6��6��gF���]��j���k��}W����t����7��+�װ��|//ܣ<�7�w-x;�[jSX"B&.'��i�^��0ɥ`C`H�K��+��꛿1Q�)�T�)��;̮��������j�B����@+�v>��ޭl^�sr ��t֕�6%�Oex̙'p낕���oH���H@�5�O��Z~������1c�p	�VC/
��G ͫ��i�N���V�m�amUQq�^&j3�S5���W���죡I(-�@ԋ�����mØ��b�&�o��$�km�L�j�v`.����ohp�����w���yЛf���y?�k�=�d�8tl�����;8H��x7"�%�1�w�`흁���@�+o}A�48s��<=%oݺ�te*~fv�{Fj���q�F���ֺz�>]��I���b��V�Kg�R��pp��Ը4I2�ۊ��Kτ���H+��S��lo.��fKP�@�KY���D��x����.�Ч�222	@M�$��)))!�'��K��7n`"��va����AO���X\�����o�|����^tA�tB0�ia�]D��?��O0�O�0�G/�W�i�?Ԕ~�u6��A�����	7Gǫ��qHuWk��gϞ���A��_���]]W��紴�a�z1�T&�«y�RS�B()�s�,ÞC��'(���7���CM�T�۽hc��0�zsuf=��x&p�J��������y�襩BuD�_r	~�;�bra�l��Q^Ӊ����-�1z���Q`��!BBB+!�Vi���3�-2�:�����Y�7In͊,II�}�Ƚ+� /�)@�6:�_N�M?��{YVV&�2	�g�&�R��4跴�C�M]]E����0�gt�7ɴ~�<^�Dډ�r�5n �	��f�j0PxG�,V�U�����j���n] �)b��.�:ߍ�6�环n�T�K#�g��F����+J\��E�\"��+��ﺃG_9�4^��m�!�8}��5��ꗿ�-%�ʍ=[m��F�u',�/�o��gH��?E�|����唰�Ie����)ur~)���\�ܖ_x!���i��3@I������۷O[��0e�_��ѕz�;y�Ѐ�:��%\1�ْ�[�Z1����d���߿��R;�^{�h���6`���	!��:�M����ޥf��k��.� �
 ���Ƹ���V�4�k���T�/6d��㌌�l�V�h����={�
K��w�����{'®K,��0{~���4��m�Vַ=��HU���I��p:{�\¤\�2�^����5�)����p�Of��G=K`���u���&��c3�i��z�x���������)�ԜX���������x��x�;�/�4����ə��l!dM[j��G^Z�fZY���YvD*�9)�ptt�=���q���|Ww�<p�^��C��ENW�j*�`2�k��:��W����(az�tkoo�p��s2�J�շ>|��0[]ۜz(��i45�_�a�r��O?,�x&��F˔.�d)��5�O�衚mvnuU�%�
�O������Ͽ2��\�tX��o^*7(��h�<__��N���NN�9�P<p��i��	_m
�n���Z[[iJth��%���oq�xs�-����R@D��ʭ�J�''��l�а#~rn��\H�g�Y�ȳ4���E�~��Q�z�z�b��V�?��G#RjW,ɂKffv�z<X����f(w����X�����ɳg������j2h����ܸ���� ��Y��������
"�ob$��ŋ������*}F��ؠSbOF�l'D��vc"oGUR\����;R��)�)By�}8�u�>@���N?~�8~��ʕ�_�s��}�?Jݸ�`�NO.��Xg�$��Ik&⼨�Џ����GMM��U/��G�9轘͠����3���yO{�P�	ooo?ꖧrI��@��ń��{i�	uʌ�4�gH�M<�P�6��/k���mN�P!��Ѷ5,�/��H��{�n�� ��k7w>fٹ��kX+ӠX��ڜ��������'(� ��9n�ݺI�n>*����c��3"�����%����k���<�<�U���y�7ׇ`��0�A�d�:�j����T�0|���p�}7�ٞ��ia_��j�������|X� o��\\\bb��;:��ii=u��k�Io,�_ xZE�{G�{0�Vt�dyx�mAb|#9�S��	�Ð�����&������Jt���O�뉎o<���	������***�Ʉ >�p����I�W���;�|
 ��'Ꙟ�,�Q��AË/�Q(r�����h�޸9�X�ܘ����C��7ɣ���VL4C�xW�k��s3ϋ$AĀѩ�Q�O�S;������� ����
L�~ǔ�8ْ �-�tWg'cC8?6��L؃����4}��HC �8��m��=����D��-�
[��k�;�c&b��%n��=�y�r��ӆXљ��þ� K��+M��+a�F�?�gRJ1DV������^o5z'>���%#c�_S�q/�?��� �#L|��F�'zd�7mשD`�����e�Ռ�G�:��K�o���N�]��1�9��u� �������@�0�;W���^���D/�X�8�6Pᙫ���vto��Ԕ�aO�%�>Uc�pu��\"S;�;�>	?7"��+�P"���8B�$}���sQ����`wm���"����Ls���)�&7�Vr-s/J���[d�ͬ�����M̏��Λ���2��R�P�L��%KK:D�8q�x������Zi�8v!E�3���ʀSp
��twW�Znq�!a?���>;�S;���Qk=�Ƀ�������s������.���zI���Z �+
�Ӗ<���l��HSn�z����h�zq��^-6���J�y�6��y J��J�{��࿒�kݳe��G`��3�m�����}~�����Ƌ"N�j�R���)���NwPc�v}���(%l�c�M�;�/kC�֢O�����ʱs�$���3��VWZRr�xc$�G�1�f:�8DȃT�jx7��װ��E*ӊ��X��7Z{�UjV{&\{W;�/�@�o0spH>�"��f@�7���?��Ӱ���i�_D�����i?��(a�H<L`�{}ȟoo���B�٪�h��cO6�6�JW���;����<ZGy��<�&l���#��R�5���Jl�}������ߔ->����AH��6)�������M.W �G��E�����j-�{�v�Pѷ566Fx� �f��_��ٔ�F�w �?�7l�V�u�B�>���1�������,n�b6S	pDdk6;!�UPP-�K����5���	|'0Ӵ-��L�
z�!�c^^&�3�� �]$l�5l<��l��L�8���~���[A�P�{�4���40���|$�
� ����]f�?�(zY$�q��8�:X�|��XOw*�!M��U?�	�lo`9f���S�����LfWs�8m��_���moo����T&�A��A/��R�f�ߖ���sS���?���?`�u�7U�GD�H�{I��C:ZT꼔w=�m�I�����O��߀�j��@� �����7 ��Ä����:�~fޠ���)Ȑ��ly�+B=~����kaL_b�$�5z�ǲ�`v�(�ʁ%�E�%���>�߿�)������B9`�H=$'������ī�4�+��^�N]`��k�]3�ք"�3e�I˱z6�šJ�KD�T��f�a�j�p��"i{+h+bu��6�rWQ2!�	_
��0��0E)U,.8׊S�s�����싱����1g���,w�O�m��mmn.-xU_���	�7�� >k�G%u��o���XY7;xH%�� X������L�a�B�������Go�^DnG��ƭIg����" J��~�=�+�Lzm@����X�k�	x^�`�hFq�m���߿�X�2e����R���rKf�"=�r��'bQ�	�,��ar�dT�I���Ϗn'EZ����>>L�
��b�\eK�Up����N��p��7�5v�//�*�&m�k�?��^�$M�%%��F�Pe��B�J< ��,��s6���2im ��w�gi]�B(�"��[���%%'��ѿ��z[�4���p��9��3a��(vH��e9ϙ�qip�z�ߠ�`�vi��0O��5޶��c��$%9���X�J2ڠv�a?Y�"o���W��v�DS���c��\�����w	���|?���0{���[]��_���,��={����lT�z_W���^�����X
n��M+�?th\��lBt܃j�(�pSKT�x�9e�)��򶝊���N����p-� j_����/ۚ�γ�*������+M�>�9 ��X2qm�� �P�G�.I���&�]]l`�	�>�Akݶz����>y8�.<��K�e������ִ?���pz��->�*]�:V9����Fa�hh�׎�
ə����æ�m �c�&�q���=��3Q�O���������i1���)%�hq�5b�"Bd���W��'*M��2iNUM�F�{�e���S�W	������Ů�A��pi4����%7�8�&'_jY��\MQ��^Ǒ_e(��8_'��ǚތ7��#���H�O���Ƭ�YWc6E�	�ٞA3]A��c���)���0;�/�&���� ���EII����@KD�^Z����~��G�MM��lV/al:'��5��u����3�Nt�p2%��E���$f`�ݝ���E��i!�'�D�{�7��9`��a����`��\��1�c#�Q*|=���J�:���ȧ0��%�:S[ *���I�c��̿���5�i��	2A5��F�C ����n�yj4m@� ��
{����lۑ���
�m�[��쪃���ے�/:R�j�HK0.�R�����' s�"��H�pϭ�+� D�5��x��i��!�$�"7�x�
K�'�M�z'��Ђ*�J2��V��\LS����U+���)dE�c:c1=Y݅vp��nWN_�O��/�J����\�[=ؚ����CQ0�M��	\vO��Anq)�w߲�Q�{QYҝ 
�;Ea��l�yef��1�S�ST/;��2������p��ZWIII�e,4��.�<��Y��2#�a���Yp�~��UTklWW�z��`��Lʦ;V��E������;�NG�f߾x �H�I��^d���<�Ԏ3�L� �V���mI
P,� Gग$�oj��Y@�H3��Ѐ�\E�R��ۯ�ʷ����/�z��������V�&���:9�;��6dMNM�ˈҨ[�W;��k������?"��)w��)Z� ��ԎM���􈾯�sj&m�?%[�����OK�m�O��$I�>�X�3]'2�?r҈b�����?�n���sK�=��PI��ƫ�Ӗ�/�D�=m�K�/���� � ����K<�7�Ʀ����u`x��:�V1wdd$�X�11=ĭs���/^��Dd���N\���G�l��u���X��oF�|�½K᨟H)s��q[�����~��)]������mP͘{�����L�O�<������q����7T]л��@��^aV�sa��:^M�/\O-M�|�!+Ly�=5����].�v��Ġڏ�Sl\?ָ�䧉�����*�-f���ao%KH�"�й�><)t�����9����{"���.]zMSI-�L�;���������5=�.G�����J
TS����?�Ί�������OL��C���-K�����[����@W� ?�r{�95��$��X��@����\_��Xox
8�y�:�>��	�{��߁�;�TUU�d��?���s�b�f�}}})֐�|Xɕ>D�~9��o�_���9�8=��1�u7M�2.c�ɟI�J:$�)4�3�~<�"��)}�z��Y>�� �A��w䎒R��	��2�?=<=i�S��'� ;S9�D�!����F~X-�����___�]��� y_�YV&��aaN�����t���|���cY�|G»�H�����_�g������.�4tu�'^��:��
���7�f�	���
�묀�P����8���Ŝ���!:n������>�����?��Ϳ�o�� ��/"B�P��u�y���6��w����� �����G������D���|����� o�o��4�h���M�h|"�X�N�o|�P�i� ��$�wƗP(����(�t�08����A�[G �<׫T���T���Ap瀌���������x��!ʠu�V|w~3�;TPP�#3� I��o��=����=d�X3ǣV��{SD���2zqf +Z/����b&`�	(,:u9 ���_��� ՠ'�����KR�
�^��;Ӂ�5t�4J��L�UT����@#c�knn���'@�����%��J��n��!B>4�%�$�e�K��^)(��0�TU�<HO��{���gPb�p:ҁ����ӳwr�	{u�ژ��Apz*0��Ƞ:����§}��k9�}�[|L��:!r�Kr�#�Wғ�|aI��+�F��D��;��o��Ä�=�!��!O9-�������C�`�-�����i0j���Y��Sl��TϬ��egS5�i0��99_8�gO��������1pv���������t�Q*=@<��+�D�f����{���1!^5�ttt�fa�к��C�(��x���v����z�_�_<2��C�)�����N�G���%*X�ly��)r�,&��K����O8%p���-!9�ؐ�JQ�昶}SNYAO'��?������&	;;0�q-�a�H���.���P$�n�<�3H#�" =�v;������G���Epnn0l�`�7�ܽ5�0V��ה����a�hg�����ŗz�lby�G��9�}���Q���@����9����ꪴ��"��^e�/N+�x{S�N5��$��?�`Z�ݸ��+�e��Y�3^E�;��d_^��dii�ՙ�/?��B��+���a�r��Jyj����d;�v��Im����e���V���P�^��ۺ��s[��wY� X����0 T?@���0��P�OO_�[_����R�T�`���5�́�2���ʍ#`�n�v��ǒ�TZY[3��+��a��%ޟ8� �.k1 ���N��)k�uy@oO#��!����gZ�&�䞵5Brj�_-_�N�����	�V<���;�f_�m +���	��R<Nd���r�h��L\\\�R���K����y8��J�5o�#0V��� �;�8*6��4����Դk�0Ε���m<n�C�*��ֿ�Q���]�1 ���>g�NAPCs���)�F�ި�ӟ�]a�>U,~�aF�+�m�ʓl�S��q<v ��P��ד��=H��ηփMx����G�l�]ӵs�ͽk�F�9�7s�
[]0C(�?	��P/�z��J�+
E~{��FCC������{�޻/o`����Ԅ΁���w�Ī����^��<�7��<��qU�#DX�����SFg���S]y��CYXY{u�T�3bu�ap��#��Ն��j$�ة�[�x������Vه�?QessӠ+]�6�UL�6�vmmo��5s���4����8��� �@�~ N�e�۫5C�E�x�]��,�<M��~K�v��"g��Q�g��U�m�_�@ʖL6D��+H���) �Πh���.�_�������$������1N��*Oᢼ�����B�RV���z���[g����h�Y�f��k��ė��Ɩ�?�-�w�X1_F`�������x }�m * Ѝd���QR�]�H5��Q���9t���g���,-5L���ݒ��
�F,�T�߹9U�Ct���z��w�f����C���4Kv^�[Z[C֒k�R8�	�`b��nnm%��k=������<��t�U����a�(����|,/�@N�-� ��\����0��#pyF����W�Æ]�l����v�!�*�/||]]E��Ow����� ��ށ����u�&TB~@1������[�|�2�`�E�C��ga�Vny?��fd��)g�G^��Y��c�m�g{��<u��Wu�� p3���6�<�� �d����Y� r]i�ê����mL�:��￶{7��}�H��7TVf��no�ȑJ�Ϊ��³��v.Ľ��â�����L$J|j��a�P���*��&��ܹ�眒�ꪨ���Dy�ڨ �Y��I+J�(0ŕ�/��s���_��^ryM������w�Bh7��}���"}��2p�����G�a���ʈ'���O� ��q4@���h��h�/�p�ŝz ������=@-�6g�Ņ�w[�����Iӕ����2���M!�د
a7��}֮b/Ө�";{^��D)sss@&�)C�'�Q�_��.����S̳4���O���H���j3��\_9�@����aC~�{�.��{EP��O������Y�1�v�
���o�'��g��"&:a�?ܵ"�k"&�yrK�k�Ʃ����c�`������X��o��Qޕ��Qt!�������Lc�Y�Y��:�=,�ʳ��9ӂo��e�ҟW.`7�QWN��� H,ಞ�{�g�Ҁ�������	
.'��	�L������ȢM���8x8!�>R��+��}��q��8���@G@V�)��"�洴4��ۭ�k@L���G[4\8!F�����W�ܶW���M�:�h�ҟx�\a��*�}u�q[�[gZ�y�_�-.�p�s1u2
��of����
�������SΝ6�{^�|���L��e/�rp Q$�闛.��a�q������ͭ. *m�QGvn�� үjq��]���t� 0WX��J�:���_<�|��/P	P��|t,|��f5ž{�޶���9Xl-��8s�(�F#����G��z��[�2hl�4���[3���p��X�筭�G��,d�T~nR� ����=.��d ���8�I�%հ����9�
眖{�j�)�����8Y~Q#��]pd�����?���ի���h��K��(uu���@�큹jٓ�����	0���P������H�rF☡k�ƞb<	z��vp����j�����J`�����ȫ6d���l����6��|�(�52u	_�j~�Wz���3$K:;;�b�d��+N���\#����CH5���!��I�jȚ����z�hƏba�����^���vM���BA���!F���;��҄ُ�92���lX4Q(� fn\栕o4���(� � �?X����_���&0����VV�NQ���?F�t��Ēݫ������� a:1ti<��r��P�3]��!:YZZ�ܶ��A�4U�������g&:(�1��{���f�������n*&fb�=GO�F�EO������a'n��AK�t��ߧ�T�-�8��L����A�x�9��,����oKw?^�����T�h�t�W�P�wW��~�����}XR�+*��m��7����Hoo]]ݐk)	Z� ��S���zN���z9.5��D];&��TW�+���^u�H�.<�ħ�2b�\*�e6��5k���w�����=^F.Y�ӣ&M�{ZYYi͚&c{H$�d��v&j�����3�KZ��62��a��������yBV�iyk�׳5���^>)�+��y#dA�g���\z�ocO�]=ؼG�ux�������6� u��ϯ#H�4�� 4��p �S'��K�n7�7ɇ����Ԡ�R�}"�N�u�[�������H f�]�, d�e�&��J�m�(��6�읜j���
�o��{ccuo���M���e���q��Ж����	/'��~�<�Ιځ<<T͊�[[#��2� �%3v�� T��g��9�? 1�	́U��D�;ڼ��R�T(��@�p'�#Me_��D��`�ޯ�X��2�y���EI��qɚ��1�L|z���������y��j��Oo���,#�P���I�䜩�?�r.���e��TNa`gW~!5����211�N��t�1bȗ��W�^e��������s.R���Bdԫ��\�}�r��>Z����/�;��TYχ7d��q s�����I�|!�,t�p� ��5�4#CC�����2GJ��ᓓnQy�񲰳oW���LȜ?� yڶC��h��"sc�Ѣ.�I��������O^�r��޼y�ݐ�����pJr�Y:�E&\TT��Ą[T쑻WgvII__Wz�L𣩲�������9���333}�W7kCN_cB�B�<֧䩔�I\�~�b�b�j�X���m�Z!;;[ t�Qz�J�F��-]]��J������Ed�~й�9Y�Y��
h���e*��:~)��zu-�f�l�[�����f%�'�c�<%���Jr�x�򝐜�c'��>���u��5F&&�h{{������@�C���0��h����9���0��e�8MO}�j�ɌH�AS˃-���^�L�tWB�/cOV]�q�<�cL|7�@P�%w���k�.-=���3v̬�{��wjjj�5.r��	�*��0�޿p�rIKRN��~�a-�Q���]yO���C[�,��N���BȨ|4��n SØ���y���2M�`K��TI�5�逸�v�;}��Z؄����#�)�,P��3`�a����9# ʗ����:��rՁ����ՉV���Oc�r�0P.q�`�wzHԋ����Jw�9w�Ruf+���9m��+Ł�"p�0=��կ.]��]�'��z���l�^:�>
�b�vq�B�c����8\�]�* =ˇ��@�5 � �Qy���\��;+''����qZ������g�r%�|��HY���>0�S��や��n�`���(�_3�e���ɳ��E�tK��k�����nW��Ĉ7T�?��� �L▃���{N�,��Ǣ������>�X�Y�)�|D!H�ri�q��~Tl4]����A�i�`�땺2z:���|��دCi^@@� SA��&�4�y� ��԰}4t��� ����f���9�)�ut>�LM�JZ�j#ȜB�>���Hm.�aL�U�Ĳ~C /o�ַ1�;Q>�W�Le��~�z{��Kψ9����2���Ӿ��XSSs>�-����q�.�!�2�d��)c�ƍ{�������i�����oS�F ��v�� s�1�/:�F$�K����Q�ElI.�>�\��u��Â��'��Ɩw�FN^#��t=Gy�F��d���*sdC����e\���	����<��������  r�3�uY����_)SG���čE�9��{QcmгҮ�ۃX|�h� P%x�x�if�Tۨmtц8D�󭜮�w����Gs_�XGo�òD����b�Z��Q��u:XGiM�����d�-�v���@��;L���a�>S��Ο�S��eC�>�-,b]����F�t�2�Tb�[��?)$����}�ڵ��PY�..�@�lfZ��y2J�)���%+�U�D��eZ�g���,��ާ����=��W>6�r? 5R�,�{p&!!����Y�	����I��z��Y�,p��,�o�u�����O{���B ʓ�QGw�/�.it�T7�����t�˰xv<4j���Wh���\I��$ly���_����N~~��F���k׽�@��
�Ǥ�;�V�@��=����J���T�^�QX�L�n�tV}n�R�c]1Χ����9��s?�> �Z0l$�5Q�қ�.PȈ0���1���ۗ���������� ���w��P|��6ёqfHJ���eC/�c����# s�7i^�\�&|x����*2�}��_����w����?6& 0&fQv��y��KH����l*]i���nT�$�j�e��ޡig���Ĥ��XsVXx�!@*�Ռ4D�<���5°������|zz��j��E�3�A�b55�;4y��<���)�_�m��4�����N|`	������߸���^�����xۉxl��\�uZv��\���2P�WV]K�#5uE+.����D?�PyEN�� �1lllb�EE����R�<������	�u��-��$�4�5��>��'+J˨����s ;�<<U-cߗk �K��9#�N��u�����`py!~/շ�vX�KT��ZG1�4�U �8b��>���BT6�HH=썝>������a��&��0�I0�r���׹>�}�W�+�ǉ�Q����G�y�.�v.�嚋Z�t�M�%4edd W�f0�)�������.�����tt�jjj�w�����q�������"���Ffb7���QK�9����s5�Kf�`��O��.�wp�ey���v����J�ͮL�Z{���`x��+++B�ղ!�I��t�e~���꫱�S%��'�R�#'��� &�6 ��X��gZ��@+&'%�k��/'�I(�T��X_Qy�����S;�j_K��%�}v^���x2�Z[��]���`Qdw�'!���p4Y�0??��H!k;כ��ճ���r���u�r*�O ��`:0�>���:�+-���ʀ_���y�&F��R=���K�V'.g/|����[��E~~�Bm��W`sNX��[ڙ �����`.�S�X��������N�-�\�Q�O��&i,��La��VSD��$Age���-��˿�!v��3\&�;��H�yɀ�N�,�θē�n����ζV�jju�|x�Z��~��)L���3Rt�;0��(Ο����Uj�CU�l���f���#�EZ�@�Hi3�����ᮦ��
f̀=׆�W?����O�%w�4��eM�jBǶ��>ݞR�4��e�p��?�@����C9E��9~�-fB�Y�(���* �X��6��y؛�D��� ċz%`0��\�7�~yt�֭C]`���^>
^����0O5+���sۤ������&Vb]�asK��/!�Ǜ�KM++��c�W���9�_�qe"nk�)/�093c��6�W�)(�>᥉u��� U�
���I(�
A�H͜6�W����3n�hV]�vp�ys%9�2(}�0��IRe��� P8��+���GKK��Mԕ:˾J�@`������	�R0�Bm�/^��!��D���,��:���}�Q�d�*ݗ	����f��d�`d�����I��0۴�f�^���Y,���z�ڛ�u�ؽɩ�c[wxF<�"�#��'�e�����R��ro��W�N����n�e}Ac"����X:�Zʡvk�mD�n3���`��>-K���c���o�����{��<��T��
���E�m�b��z��1�gSwT�=�݀���n���p]�zL����Va�bXN)F��"P��H��aaa�f<� qr��^d��n����1Szz�ܚ%&��˜H9c���_m�Lu��k>`r�����S�y�=errv�����:���~�P;^�1_;�W3��}��A�$���q�`��|��B�8���1��;���c�RA��ݐrv0=,zZZneC�,Oj��n���W,�?WY/��5Kh�yZ�p=�9�s��n��P���^w>u�؎}-���E��6B����g|by[�&0�~���*�M]���ϟ_p�xR8>� KG�,EE��o����!�1-�N�MF�W��z�\���<08�BL@�}m�o��rZMt~˦&C������d�z�1j����c�tE._>Z۶\Ξ	��9'VVV�&Eθ+��������Gp��\�!}Y�%����1.�؟�,�uh���"�������!�W �]pW���G�@�"��_E���T 5�Tf�M�2�m�"|��MBBf3��!�-��r�c�������ѿ�@�u��C��<�%ܲG�m�����3���V	(p}���N@����%��Ux�+����d���eU�Xa��A�U����L1�b\�ϟ��*�u�X"��{�'Ⱦ<=%���.���л��,��8�6����rO2���{N����8��� ?Vr]۞���.��q���م����&t8�����e6_0��X��t����H���`/���~`y��j#q��������
�s�qV�N#���2��Z�qWN����W�_]���'�i��<�;�����:I]M|����T9/��V�����<w^�1)������-�������.m�x����\�F�������1��$�ۑZ?����M�i�a��o�wu��3�UUu�R儑��׊ʶ��g�7��$�,���}bw
m_K�2�傛O&30$W�2�l�Ł�e4�ݻw&/~Nϔ~ڇ���<��������.OT!9��d(��

f!����B,�W2R�~#����`2�H��}���G�W���V�8~��Љ�V���Ȩ}v�⎂�t�&]\./Pְf]�𮪞lcx���FY�����x*�i�懤t44|?���[�{B�4�[�.��ÊeCV��FN�::�ɣF��㥥��*�����֞�%��7�!"NO�^�smN]|GGwx�JH�|��V^�Q1.漨%����p>7����>?�BE����+��#2h�=+��_��ŏ�.`Ǟp��`I�������H w��K!��j������7��~���Z��d����z3�j�.�� ��;�X�,<�VR*�JH����D�\�#O\qB�?�1q������{]�*C(]B����5]����DD�Ǣ<����o�	a��=ɱ�������;Ew;�/)�Eԉ}�1Bze�n�+R��Vr�|W.]:엪����:���
1���s�M79����7]<{�d�����%��y����ϵU���홊qB2�ѳvX�uj��\v�Z�%/U���U��յ����~�'���*ӷ��el���z0Q��P��P�`�u܃�ϟ��-j��Ad PΘ��nb�o~�lH�9Q��*��'�����~}>.�FG���8YI���m� -]��v���2��"3Q�{����ApTn�C(�C���=^�#�Ew,�ްAf7D�=���UuMM��<O�X� �w�� ��ldo��d�ۛ!ܩ�j*Mu�\r�0qւ�MϢ���i��i�y{�g�'�k��=*;`Y�\�dA�
��a�����JQ26 ��tp<��u����^�,�5R'gF�L7L�*���P#^
W��^�	Oȁy��!��sJ�~߆*[��M�c#����Ѽ��H������)F��R���X\��h�.-=�`�����g��©l&��cq����ι��wCN����\p	`����r\��dF��f�h��&v%Ð�Ǹ2x3l�J����,g����TdtEn  v��[944T7�ώ�I�qS;v�Py�FFZ���>D��#Zcw
�Y1����+~���3H��������E�s���Y��G�e�Z+A�0�V��C��DK��\�u8�懄r|�"L���4Dk��l;n��1uLK������29�Z�z��P�0����hW�R&��������d��������ͣ�X�L�n���5,c�e�����E!�R~ڥ(�c(G��ܵi��bA���`����;�����߿�?��<����Rt�h!R!mHDBL�}J�%�RJh,Y�:�[�P��"�����lI�$	1$�g�n��:�Q��������}s��u��\�^�l���J�����/B�|\(@����TպOoP PW�Zv�J��ԛ?�7;#E�PQ�HĪҾaΗ��������V�FG㦟�����t�q+��/{�#�+�G<�3��6r�;����)Tc��G��Clk�������Z54<��;W���6p�}��]��Gx�\�I3�%��X��x�m�dpr���z�{�<�?ix�)����y�/Y�V�
��o�ж��;|�9�3W���p�!Xj�J�:J��p*�1���|ϠK,v�z1����T�8pO�y��K0D2]��^^O���;�c�z��G��W���ǸL�Е���_E�pKgg�'��m3$?H#"Q� �o�uk
�qR�q���ۘ��_�^��z·Lan���y�P��@Z5t�{b�O�7=n�)K�ڤ�`^G�C��$�c;�Kz5j(��_`�>^H�K�����3S��!�=`���잼�dԗ�	J�p��6�o��ۀ6�R?V-��^yy4>:���M�ۑ��-乬�]�gmIi)����j-���a��z�>ze̵�B�?o��W�H�?�S����B؀�)Oj��7��y��1�m����=Y�$ʴ��t�^��S���0=�D'H��vo�X �N���
�L�ZK�*�=������&�q_P��ЖSV;������F�J)?�'F��F�F�H2�e��}�P���i+�~�iq~�s��$�i��I����/{�|�z+{v�.��9���D8*�g�7n�8�D���2�gV$�G�mܗ�W��b5�V,����Q�Ý6�&�
��@�at��$��ǰ����?�SWS�{}�P_��ͥg�ζ�^��/��)��9�����}?~��~_��5j� 'g	b���'���?:G��l6808TR
�NS$��5}F^��ȿp~�^���e���9�S�g����Ǐ+L���� x�7�K6B�Jڵkz�]�h��}_=~KJ\ڒ�-/���w���}����U]O�?0�º��BM��x��TU�b��=���en�{hs�@�V�Xq�C/M��R��un$�}�|�
rrryϟ���F���J\A�[N���m/H�Ukߔ�����c��8�d���r@�R�{̹�>C�u�� �L���&��56��M.��A��=����L��""��T�b����+Z�CCS����*sR��p��ay7Cq:���.3����U(;}ۃ.W{������ꪪ��:�V�g��6���*'XҜ������t�l��$�&PD���ڥ��UXH��������{��WJk��}]��{bov_z%�4��/k(��K��v�`�b����nO��I�G��͓-���a��Y�粬,R߷�v�%^�2Z<�-���:2}�����nuk�̡3��w+@���6`M�B�l�����p��^^�).�������9p�OH��G�#3%����	Gŵij�>m�W�����_��*;K��رV���KvRqC'p�(q٫����	�\�mj,��P#����u����]�V��M�6���W�^�%e7��F>��.��KV_|�+�'@&m6L*��H �;~�����##��x�Ve�����;[���S�V��/Y��aG	®�5�5�)�F��25�E�� ��$��bwd��~��p|]��]	��2�ک���vm�U���_̯�����V&($��In�qyq�\cS�%.���a�J3�$8b��!.�����<p퇸
n����]z^Ť�+�j������&��V1FZe�e+�0Ni��m۶�!���ͥ��VY���:��T�����s�����ޅN`�Ri-�5X!�q5��C �]�ڀZ��7n����2�^�l9��`�Z��MWՁ�Pv�;�3#�ѱnK/����юϧ�>Tz�{�ҍ���O�~#�o}��.s_���,��(e�J���	���j����k�|��ϝ�X*�p��f3����x���0�B^B� �m��K��|�rZ�t��44�<ILTǶt����Y'��ή{|U��Pm4��͏�8XBSi�ﰙ�m�^�˯���*�;���-Z�ĝ�7��^p0�H;�wl%��]}�^�IJ�>ܳ�y7)���F᪞��1;���@���ѐu�b���өU���������|� sG�����x^���<'�ԕs�U\���,����HK=,�� �$׶�v�<{�gT[UU�5� HN�/�	�"���?z}���q�Q�K&���O�h 1��/{�zǲ��\��˫��:t��a�~���!���O$���H9"o���}ժU�i�!/��n�i��� k�k�X�HH�3��H�c�,�Q��J��W�u���Q��4�Zv]��!��L��<�*�V!��=��$�"wY�$J��is��6���w�r8�-�t�^�rt�x4�,�/�i�O˫�?ތ�J�u�Jج��Ӻ(T���/��^������ݹ����.'�LO�=u.&c�w�Vl��;�woč7�&���ci/��V�[2o1��������DB���`�;�a'�F>C.��]�L��Ƞ�?;N2�V"L�AF��?�^��?�8�c6'cKP� h^�jf�����<���ߡ
9}T�����]�O]���ksp�Ӎs>č\+��\��$��FL��M�t��CX��!�!�����g�0�J.�5uu+��$�G��"��l�.T�E�����ruq�9ZY���0��~��Y�r��z��$s���5��)�f�>�E���1>\
� F�g�[X�u����\JIs��ק��#���[yp����S�O����_2�(9���X?�Y���K(�����m8��� �~4}�=���븝������U(	Uރ��_8ea\�n������6��s���zBs}�:wNa��j�)�C	�vHM��M{��puiH��|��Y��-�qbA|�̑֎���pDs��X���e�t�[::ʂ`?a�ܼuM	�%�o���P��>�Al�D�P�~�#�=H�ҋ(�_�7K�g�Q�bo�O�Ku�^Xy[&�|�Qq-��#���%���g�d�K��\j		56?JH -�qVq�U%�d}��8
��uU�dnI#
�^ן��/��_>\�SHe�b��Nd$zK	X ]��,4))I�k���Y��чh���f��W���K�ݏ�(��t���;����9T^���\�6���YJ�?� APU$'GY �\GFݻ(z��\���]����~7B_����f?�U��]l�{U���I�o�t,	\�n�-�Egq�)��]�+'�^_��0�]�
�r5�����ɖRi�+�`G��~>��a~MI`����S��������@�����3�(	����]��J�����;�^�|����G�ݦ�s��4�p��ى�0�-�M�K�R���7լ�,�S�|��Y�U���{j+@��vvj�2��N�ԥm���@�@\Cg�K���b�Hy�ϕ[۸�B��_��Iy�"I�{c��fs-MM����M6O<9@�2J(d!�o[�7��k�Y�� t�m��R�O�	5�c����{��������X����l?nm-��ŋ�wk@�����S97t��b�%�5��qj���p�`�/�t�s���2�p	�;�pMN�R,ok9;>T��0�n<b����>)f��2�$��9_a���࿢����/Ꝛ�Xp���\�v�kܥ�n�������U��|��;u���mh_�V�(_�[TA��k.͎m�>�hk�}=<x��C�IF^A�q�$#���5�FY|���(�d��k(]흝��T��,�(��Et;��	tq����[�`���gii�8/�I-�O1��דb��e�=���Û��[Kq ��U�yr8p�g�����m�M�Z8� �L�/v+&����	�RL{.>}�A�5�nKc�����'���ɱd��J�L�gsfD��W��+�Uܜm�wC������@̈���T[���W.:�u%��~�ytM�>m�̭�;C6��y"}� ���]��W�X�����v�ɉ��ć�Ss����G�~mk3��No�����"���@�LTu8��TwBN�8���
6y_������ޝ�����gSSC��΀@�N��,4�4浝�i�Y�Q)� �ujw-��9W-���d��R]]}Dj�4K?=�:9Z�u2��\���Hw�[�V�c5���gƉ�w�/F��Ͽ�5��Tg�����c�n>a��;��FN�[�_�b���vkLmW��<��&D�|?7GZ�n��c�`A�����M���4g��Z�����!�^z��"�9�q�up��9�]�\ʷK��C8��}<˄��٫�0��~�w����4��BA���7�M�&É�^�K��jb׭~X�����k��yn^��2���	N#�\����w����##JD{{x.����h4���էW^�T�_{a�p���}���z�4n�Mط�}�G�;�����&4=�R��:��� �HQ��o2��x�^��Z^�9a������kN���1���b��[�s���}���8��%��nr�z8��"��/N�H4�|��d'�3`��K�Tc/����0'}t�("�'q t���>2�éRgѻ��{�'w!����}H="���-�n�vF�t_}���s�=���A/-t|T����{{a��
k��l��{|N��ͥ%Qb�Z���ck�n��2=��1e˷oEX���]q�^���&��;z?)�E
X��Ees#qxUB���6�-�����b�#�M}l�]�^gg���<A/EEt4��"�9W�msZ	i�1t���Ϟ�;3?��A׋>��^I��'No���ߍ��g]\�7m�$u��k@{�-}�����w`�5��?X�R��B]P��(]�	�
�}��C�WI�5O���ȚoZ����j��S��Se��JW�Ǉ���d1>�E�h��5k��\)m�Oo2ى�-m�Y��aa�{}CJ4����*'������S���/��{i���C^��ZޒL�Ϲ�6��v���7_N8�pdyk�Ÿr:��F,{>�a�~��ל�yn�8=�?#k)�rxx-4w�g�@A/��oqd�������Gݣɞ�_����vw��U��B��ӣ�:�DDD8��$��5�<6H��B�<Zµ����pB��ϟ�Tw�N���B���\����j�}�Y&�A�Q쳆"��7�f�[8�y	gQ���k�@A1H+��Xt]��Wt>0���ߞL�3��F�.#A���_-,��*����\�k�&ff%�����؃�ܖV   ��,0��5����єۯ�[~$�]uG�А+dud5�C�Pzr���2��	�k�˴ؒV�;w��}jI�8���,Y �2�(���"Dz:��'���n��6>>>�F~�W%�����м��agkK{ПI�TRQ	��7�셟r�M7n���l�I�T��N�W�YRz��YUH)9ӘI�� _UV8*����f���/BCC�\h����=*�����X~4�D�=���
/�������t�\0���|�d6kγ9P -F3[�4��M����:B������r�~�n�F�� ��b�d����`}���O|%h���K\8���Kֶ�����}���9"%fU��P��-����W��D�M�XcM�W��'�T?��]�]@1N ¯ V^H6H�s5��Z_��6a�dī�I(�C`vz%�����|�U[��.���g�1<�����>����ظ�W���sB���`��G����B�0�usF�G����7Yi&����(� �x{��c�WMey�BAPY���Zɣ0������Y!�)��9N��s��&� OE�S۱�$*F~Ć���)�"P�m���ύ3|v���x6�Y>��:��*LP��Xݦ��9~�־j#����ϟo�L�4�R�J���O��̬���G�R �P��==Upz)G�,�
g}��$�*EآK�	�����H6('cߩ.//���eXC�#--1&��]���.�_��{}\�N�сg�_�b��!���u8)O����Oâ�14� d�M�| �-wo��g�ӹ�����ٻ�|~V��`��'����hiM�q��}y��h�Tc��h�-،��������,��(?,吸]�.+�m��2aG@���E���ک�¾�-4-���'C��ck� �XH�[��>L��|p�e/�G�7�|ܲ�RT
�:�z��"����Afy	A F����ɻ�>J9id�5�-S�ut��9�`����uJ��>6N� *�0�\zNƒ�Χ�R�<�]X�҈�Pu;L5Zq�n	m�Pā�G����c�[�*q�_獫�F7�#e�G�1��H�����ʣ�^ur���5?���~�R��ɢ��<�N/���N5�P�%!FS�΃T��w��uVŪΖ(^����z\��	�;�vnЏ;���B6i�g]����`0bx��dd��Tߣ�CT���Ł.��O�cjz;0����g��<ůS�Q�U�zٍ�'�V�Irs�O��O��)��M�<<H�RU�{$]D���Qx�:���]�)��o+����������4�,X%�8 X���X��	��;�P�$���/����>�JDI+�+��\=v����V�̉�?V�~���'�9�*h^����9zz& ��n��tuu�C@_��A���	�3���mPڢ��]�3����@�f�#��(Q�yݔ�>���ƷvDlA>O�M��nH,
߆R�<� �"d`DB[V�H����:bS����o~�9x���?��E7 )�� ��['&&�O�����0�u*&�c;O���Vw(���bv(==J���ڬ��B�}�ne���0`xAnNв�\��sn�~��IA�ʫ���e%0�ٖ�,�	4�]���>K�Ҧ��I�#u�'�����b���ވxvW@v�*�B@ވ�%�Fn�I/mFW�&p':Z#����0�-��޽{��:qll�͍�-!޲#���{L�����	RZ����9#�	��ܙ=5�Ld�~�Tc���j8(^��{��6I7޲���d�q@yM@_��H8Q!���a�v� ���g؏���駠�,�����,�k�y=��\P�C4
v���dd�+~��0��	y�q{G��w��0����-�0Y[��/�*創nW%)�8:9�]�N������w��0a���IF}:�?Wt���<���#�~8+#]��E��|���N�~k?sWt;��&|�R�N�	33��x�'>E��Ŋ��ɇz�9moia�h��wywBΝ����������=:b� ��)���^|~\���,�{h�y���f:d�_B�Hrt"�Eh�z`�O��~[o�tpHH+�$B>��r�7�r܏��?������$�B���N�D���.�\[��F�
GX��������=q5X�%*�- �5�z,sV�r���Wk�n��VkƍS��R؝Q�(���I�jyU7���J�@K��"����SA�WY�M̷A�u�c� ��G���,�y�|�D���>^�^ܲ����*}��~EPt�¥�c�7��1����������8�@ȓ�RLHЗ$g3��Dx
%5`��>��U�� Q8G��qUA�&�]}��V���ĸw�e��#���F��f72݌�U�چ��#�l���ꌀ�1}�;��Ab�!�_2N\upX���ۧp�]O1�d9������C��P¬ O�ً�R8����"4ۊ�۾���0Z����6Z��i�X�8�����J_��������.~?U0��!�?j�O++�&��N�A,��\3^ߏMMM�:� ��9[_@���_�ۣ�AL�Ӎ��|>��.�('&�[.��Zz#�t�
6O�&7� �|΂1"# ����5i�J�,���֙�yP�!D�D�o�XW�
No��8,`��C�H'u;��~�!�W���=�Xb�0Z���nc��Q9�:�t��T���sg�Լ��u��i&n,����7����[�,8\��d^�_�x�D���7�<�f���g��?K�ɕ��v�T�A�N�`�wԋ�`�X�Ӣ�~����_9)_��]�kw�rOj�{���"٫<h�?_���̛��G����(�Ì��Y��[�z�I�y"�I�1������zЍml����Tcfv6�;)�CC1z����w��V�-61y�����ދ�~��t�� m���)N��?=�E5�	�'�L���LX]G4.��L�D���Iga��0l�SbFv�c�s4���t%��lb��ꊩ ��~5O*G�����|�]���8�ul�,�]>n�-�PБ���꺂�C�ǳ��(�;�7�C55���D9��<W
�N�=j��<�d�������C��&r��M6�����c��g�^��1��|vg�ܘ�b|��x��c��+e'�=bcX�荹�u�f����<	�"�#�WЕ�����E� Fh��6w�"��u蜽|����3��}�4E�k_�&�]�"��
U4H�K�>�J���R ���l%򡿳&An��0`M)z[|��s�Z^�2	�t�Ć��=����S��i��8�&7���8p����r�F��� �''���[?���S���ʷB�����WQA��!$M
}{G��j=6=���\-��������`w�~��g�`
�K�b�� ��~��hw)���$�j:8;?�&��k�sv0���g%���[J��G�i�?`W�U555�^��X��eǔe�$Y������5�i��ʁ̜�+iiiN��&��UN��4�����S�Wd��q;�M:�����z���ς<ߴi��ٳ�~A=�����|H~��_mԈ�fi�d�q���p+"x�G.���m�!��j���!>ׅp��瓵���}2�R���N-j���_�2������z8��>MD����d�SքY�v�E����z��׈�B���U�KG�8�5��#+P��K5d*$�0}HX�Y��'��(�"��o�<'�,�?����G���j'�F�p=�;��t�ž|����J��oϤ�²����V�������x_ͷ4q�b>ko�GH���R4N4�B�2	o�C~_}A�q�pE�Myi`[��L�L���cY~��ݑZ�����ê��0n�_��^��Pw��������:��tܫ�h�B �	�a�O��B4ִ�����<�|\���EZ�4�S~��*�z�i��5�n,���P#|�	���s��<�yÏp	�~�;}�`|U�`���ɤ�ө��>����˷eE`�賍{ ���]��NH>�ߔ�d�%�Mb��U��JZ�eW�SU�a�	;{�:U���j�l!�aK^Z}�+k/���}d�aa� 0���	��Ϣ�:Zɵ�U�|���O>nUe�^�w�>�)bi���_G�ؤ;������<�""�mkh�Nn� 3�����zI���7VSN��P��~�R�~�Nl���6��C�|k5����iH\�h�N��o�^f��w�$q�U{o��H��({�z�V��N�Z�j���a�M�kV���	�"?7�����S{h���������(�F�Y�A�A�=F���7�e���-K�-Ԇ���0�x��Uˬ�*g���>+ӇWY����
�oq�T��SH�*�?�G���>J�w?L[��T���Q�FC,m�dj_ ��؞��r�!s��K_}T� ^�y�v.RCU�K�Üӗ7N<��(�e�<���ZH���y���o9*O����5K.e2}>�\?�v;`�=�t7�k�$`@nʬ�M^,,,L>_=�&5�Κ=�s�K��^��%0{�烷��gmlK��#Hx(�ɺ�|�`'����ʁ�-�d��K�% V��W��[%H�i���@����{5);;[���Z���'�C���΀� W�9s�K�W����͊�m�KQ�n��璓���ض��a� ]ް���^�A�բy��>�`M�gB<�`�Zj��\�T�tu�T~*w��!�aD����}@�S�ԉ3��KĠ����?i$����xbNa��н+����� O��/��j�jI�q"��� �@�h�7��,3e����J�ֆ���E�Ģ�k��c���=5sl�-��0��A����7ա#�[\�~�mX�IC���0u�V�W�,/�r�� �v����v�C�ѻ���_}\vB��*�~?)��q #4j���$������e�_�v�ɕ"��s�@$C�6�932��,��� ~\�"���?��722RIU5�N�Cow�Gn4+`�.�eddp��B�<�����_� '2��ȏ'��L7f$���Y��D�ub/-#d�G�/t�J)�do]]�eÛzL�tq����A�^��7���s����M=�^��J>58Y30��#������iYu��P��`�
�^�;�h�X�d���˟{��$�)�������%���r��hl3�S�P�?��������bm�k_�m}�
y��ԋ<U��2�����
�����>Vx�I�d�FA[v%Xwa:���@����8��`�)�l�c�w"����|�G�^�|�B���F9�IX[�eɂ顯�C��4O�u�t!��N��"����M����^Li�,�b��n$������T��>��@�B<.��{�v{Î�%���ӣ
�W��}�_�H?Ⱦ��T��Kv#9�D:?ª.�r�lh��+/��������<I��u2J�HuDŔ���c��8�>�TO�%�ϰ�������������gi��Sה��b��������c$_}��z�.+�����o�ڦ����oa���f���Ŵ� R��������;{4�T�@X�~�O�GP��-�H�@}P+sP���׷���J��O��K��L��0��Ae�b`��<����ڲ�>�=d9��<�U�}V.B�#nŸ7�6�hd���m���p�Ć�G�,�<s�Fl�)�}T>��	,nQ1
����fN�Y L�z��k B�p��O�ڵ��-���dZ|�Uy����>h��y�j`����|�r��%/~"�u�>�a�6�/�o;��~�FR���J��ꈀ����ʛ&ϭS��/���_�+�z�zdI�=r�c�~,�O�G�T�VR�W��6Er�|�v�	g��2:�C��&D&=ќ�ZKCZ����D��� \ њ��A�d^���
&i���ݷ�P�x���89}���*>�s�И�غ�=z��9��α���B��B?^���"=�G�G���'�n���F �s�x��T�цK)P@�к	5��VH��m�T� /�����gВꀋ?Eo~y^�˗m����n���j� �0< �I'y}�󦻿�����f������>��22,ٜ��o�"���D�!��O]��JPElk�D�	���4�V��!�9:����RGa�Zk��o߾=�������,�'���"���J��=U��~_��z�bz�F-���N�xS�{��`��PO�Y�+���wtbS��[�F�bIk��P����_�t��մ?���� ~�e����S��)ri�h����q�bٜPݱ�_ZL�Z���	�9wp��łx�������Ͳ�~��!�(�j�m�#!���	*���F6�#\<\@-�n�z��c	1Z!u+�l\���1BoE�驶
���=v¯17蒚����]�r���d/l�\����)��r����h~������<W"T��q����9ޜ�5+�S�8��ʐ�C���.����b����Y�*9� A��$֑���V���>�1Deۄ	Ӥ/���������=-`���p8��rst\:0��&��p?OR���u�m��λ�>:�G"˜��r+<�m[�VG�4�ׄ�C@"%<����~�W���FR	Y=�*@��`NtN��T�ϟ?���g2G�9��]�M'~h���l�V����"��E�� �������B��|�&��T���c�v���K�L� �:{��~h3�g0��p�d22sr��s�ZT$ň�%�Tw�S��,7�Z'�� }q/�:�}��ꪲ�YyMO��P�Y��L��!��_��u��N�9A�Q��KN�$Lg�I�Y�p��K����2-�8���=�
�š��c�֮Q_�U�0$�X�C�Qɛ+���|$`�؛%��V�����o�%�j��P�د�ǠTA�ڑQ/a �7O2C����:DA"@��O*G)���;�N<A<uܙ86�ik�2�1X�)�훺�R��c�V���;wV��t�˗ϧ郦��i��%����9�%��N��z":m�n�^������>�pe��,�1H����D?�~��kDD�,��xF��-~倿�� ��7�0�	}�W1���;$_`�8U/�W4b1��Ǉ��������!EZ�О�^�F Hԅ}p.�1�C�4��FVl�>��� A<��H)	��P?�*�w�ϰw���.��P�9�}�P�z����aMmmmk���ļ@�D�ӛ�h�*Tw�ho����?cPr�A%�p�i���_�m�݅:� ��C�Pf�Ṿ�L����2��R�w�R�[V�ܝ����}������{�4o�3�_��0����~��<#f����G��5�]@A��I�P�~���}�`<9����1�yٌQ
t�X���pjKM&�����\�į9;�M"�7�f��PI���v7z��i��t]Ͽ���	�me$D%y�������
}���W��s�{y�$����<1K����5/HK��Ϋ��ʃ_�r��ϛ4�9� ��%��
��4`4�����׿I��=U��Q�K�#�}�R�L����2ӟ1L���oLg�AB$L#1�m���V���q	_�IY�� a4��"g�EI/�,�7�	�c��#����@P��d K�Ro��|�o��LX0c�fk���sc#�Ӄ/�F�MR}�0��G�vɔ�Q�^8�����͠̖rZ�,\z�/����v��^��(����s\��:�t��!�0�S\f��P+}�)G�it;:��e���nUe���x�̍fރ5��+�.��������,ib���g��y��.�a����yO!k��~����}��a=ή%>J�j��(�0�ӣD��f�g�:�8f��d�TH��Bu���nv���0���ܒ�~��o$g�%�G�e͜L��nt��G.L$DZ��@�����۳sP�j��_�*n���ΆA�y+f�QPe�h �Z��_�-��'��n��z�*Ū� �:kH.�f����,�Y���7_g���)�������j�B^~6�A�%+���+>%��_ڤ+ϣ*F����,*:ڧ�k�'�y݌_���朻�K�-b��Z���� eC��Y.i��ݮِ���Y6T�9���Ꮱ��S����������3�x����Ɔ�y��0��%��=\�K���6�q?g��3J�50�>g�t�$ ~9Fw�l������MqƳ���e��K~�qFn)ݤ�u�}Ʌ��� V6�.�-Sڹ�Q���s`6��V8��b���Q�p���-���eGSٸ�װ�Y�1�3���%a؋��ٍ<���W��_W9 �v2�=3v��ӻaY������2��:;�S�ܙ��	�k^�p��6��r�Mz@���t�j	t?_&@�B(�	o7��lA�[���~q[���F�d�ө���@�����lp&]�C寕g��u*USu�n����n)pӱ�Uh��{$���>�`|b�<��Y����kI 0�ա�A�5V�3�J�_�,���6�2��k��l0ˣ�B!9U50B^�!��XP_��D�P��˯
9���C7iK0N�2N�k��PO�1_I�3��K�	)����Lm�8>G���g�[vc�����j
ց\Ồ,������<����d�W�g]�WP]�ߙ#�a��j�i�Y���W���Ml�7wa+���M�6U� �;��'[v��3�1/��#6c���a1M}"���m$
�������V�:x��8�|�H<�Y�G�#��ݙc�S;gH^(��v�IHȳ:����(+�̓�4��2�}�{�@`1��V>����V'�v;(q���w솩��xaM���_�Bl� � L�®_����ƈ8<L��SAv2�]l�9&�})���A��c�0��όo�'b�=���ï� ;�/�O��w!�����	�Q�|���r)�p����� KN4�.����.��l?�`3�J�:�RH�(83>p"�ե�dHYLQ���E�9�5K��ߪ#!  �v{A����:��kf,��ǻ���P ����,�Qq�T B��zE͕�����B��D.�K�(���נ�3$��2��K�J�W;l�y��d�Yrl7K�ˣ&��B޾����.{�x�3��s��ə]���[K�(,�j�X�m�]ȫy�`�LO�>�v6�N�	 4�ĽBg�4	�v@�`�F������`�
����7�o�T���W�"8g28ۭ�S_c�p��=��r�o�b���q�Od��X���B�h*��sP8J{a����l��QTe��Kz$`u]��͎�a��@!@�����	�UH����i�j$F������Cus
`�����޾��}�yd7�Σvz��˜��@�#a��xg#����1/�/l��G	w9+��z%�2��%�����j�{aN����:s6���Q> w��W�n�tc����ۿ��|�r����c� �P��t@^+p��J����ezZ���l0�h���R=�A�2�� x�);PB�+d�4χ{��E���L���47��N�%����W� ��X�*Q���r����k���	>�3ƀz�Fa(�{���%�BѬK7Nܵ$����yȗ��9����>��g��"�Y�z�Ug��E�]��5esb[P��P��j_�����cK���ՀA�ǁv_:�&��,��>�,��~�/��[:�İ�M%i�:�sg 6O�r�I��iR�,�lr ���	&���7V1s"S	�I%ע.LZ�n�/+D���#����T��_�8��L�������4
�F=z'�������I&f�}%�@zR�oޙx��c�����m$����2	=���a�%�����b��!�F�Uq|�[����,����Ä���|��n��v
wm���,!U"�����zkf�3��6��A.����3���}`�ߤKҲU���YrM�s6W����M9
���<,�:��*c�e�!=R!�ΰ0~��1G�gy��F"j;]��y|2�H@�U�  [t��A�y�����LxJ�Qf�NH�	rsBt9X�s2�H���+�֜�Lt��!'�B�_X�k� Q�[�ogVN�Hz���\0��k�s����`�!!�D�IK�{�����������U��NTT�/,U����������i�[9���{�����f 3~{��Faҵ �sק���a>�f��_�����T�hbI�f'��q6�8g=<�4������]���8�L��n0��<�݂�����+@|��[f�	�9�؂&�=��Ԥ�%#�s2���Kn?�(!8��18��j�ڐl���yX����ؚ�{�a=��w^�vS���~�=����5b��И<�) s�W��6pC#y*�������']�#��b��[��?L�h"��
�\���˯�ُ�o�E艫���_�����tD�)1d�0��$)꒢�o|if�Q����,��U@D[_#� q!�ك%�� 3[ϓ�7�y�}�|{�X��V	#|P}�l��K>�D��G34���Ӷ�
���i%⊬�9����������d�3�%��5�o<�������[��ㅳ� #�`Nȍ���!3�>�>������1�n\
jG��~x"�����>�N`f�2�5c��cC�gm �)�r���F/}�����$��zCDf���x�����P�<��(�V׵�Դ����¤0�m�-����5�b睯_]\�����\B����2�1�:F?�P��A��,�a��X�ph��Z��w*}�Y��+Ajp���b�+j���>S���K^(��<�������z��1�
蒾F �c������ 6\�� ������3�Q_+&�im�u*S���@�{���Ֆ3
_ٌ �����4�K8s�Jc5C,�5�v���r�ΞUz���O�ϨW.՞��&&nr�b��s�G�+�G��e�q�+tI>��� �\W$A�yHX$Uw���Ɖ��I�DI�2J;��Q�����meϽV���M�\�W4+ÆZ֙�f�%��o��43���ܘ�@�j�a�0�u� ���z.~]󆡙{�M�}_H�Ȍ�
��LLM����V�k���J:ZK��g"Oys�=ybt��ͻ8����1֕VEQny'�5f�d�tI-0��'�4, ִ�
��l��)[]�+�sC��*oĿ��14g|�9�g�,sa�)봺"HϺ,��;Iw759kl�����7����p�S[�`��� B�U�/�(j��ɋ� �g>��g�/�v���9�A��x#i�ݰ���0�2�ߴ�▚;�r��*�����g�?�?�s7�S�3��?/矷I�����۔קlb�����/������{[�Su��#��6��E�%�4��q}t��5"��iVN�I��4:X�k���,�C�LB�1}�:Lg֪�u���N !V'����.�}è��}`-G+����B�i�צ&�����c�n����	���\�Ӄ$�x�X'd�ꓮ@��#�^��s�9�1���픙�S砄_�{k���\r19[n���c���J$r�S��+�h:��LG��7�J��EdW'z���	�q]�b(M	�m��H{vSC>���e�H�S�L���n�J)E�)�N ��㯜V��~���Wkw'��U���˾ZoL���D�+��D/�56�7�xq�>}��v��+�k ��75R�g���ԃ�g,R
�)��a(���F^�
� �@�%��;���ё~-F�玞y��7�QA&H��,�ͧ���TU� ��Et����g�q��7��$����!� r4M���Vm�V��U�ytt�/0f�H�?��}ߌ1|�h�_��";[Dr�)����?��5� ���6�Z��23�VG7��Z�;:C�d`5�96�L$cz�?#*F.C��?���m�b��_cð�� �w�����~[�)_��@�	1� MA���:��/�]L�8ySo����)�޿�W�.UN���-�޾��S�5���QV�&�"��PEwD�7큵��ۇJ=f���klԣ۫�d�&�d��GFF>�v"R���c���g�~U���vm���_g���:����=%�Ȋ���OfWRS_����XJ�14^Cd/���q7��+�
��j�a������j`���V^�/��)����'8�t�����"f��a�cT`��	�DCCC?q��kG���В(i�L�:+3��cfZ3��u�rK����R;�����������
��W���8|�M�?U�Y�6T�=S9��W_�CՐ|�?g�t�tO�oͨ�6R�_$�@�|�|�T�%&zZ���Ł=�@o__l��޵쉀������`�I�����,ж7�����D��49t�{� ��B1 �1���i�*�=�)$�=�3�,%\����{<����MG.D_�O5�P���a�j�͚oU�H�`�d�[ͻ���IS)OE�|h���e�꾾w��}Õ�3�-wS�!n��}�\��W�b�j(Dx'�y%��L���X3Gf�Ю�A�E�n^���^�s�o���v��<������-�"0��b� b�>#��ٮ5�e���<@�A����L��Zs�-�#��%���U������OIĕΒ�z�.������ڃ����ptq���)U�
L�����ty�h#q8���|�@j�4���C�k��O�
� ����J�6'lch}O�)yn�R��4�$��v�9���6�L��B-�:����p�擰���7 9���O��0�1�F�Z��g��#�˧��xR���+�1���0_�&��$2y2�1�m��&f o�2l�yc����0	w�و��}����i���C�����n*Ձ��+%��􍳞�-IH��|�agw�:��τ��ę�#�����h����1��4bo6����0m���+QN饐�g�f�}�/����E�2�������}g�����PL�do2y�l�ɪn-����s�MW�KC�H�}��t���fA�&��V�`#c�~�8IV3`�i��^�`��k��ln��;��s<�:v,P�5�tV�8��Z~���d��Já҈��n>��� g���]�x�b M)�B�+P���TT"&t��$�f��t�V.��}e�r�_}鯊6�PRQQi�)%��� �U��b2fZ_t2��ĲF�".��d��Q/�I���g`S��[~qR�̳'}��q�H7Ed�2�X��>�n��w����ע���rch���]J����U3�P� ��V�0G�g���IG��
i���yW�IE�C��1G�{g�΋�����4
�:�\��[�@����m�h>������ˋ�s߹ ����T9O9�Ԣɔ>ҠV��jjȯ�e&����ڝ���cu��\���)��Ar��E��Ҏ���S���}��1��w�(�OĪ�u��E��Mh�����aU�L\�,��7�
R�W��{�);=�OH��e�#�'���Z�z�y&S�����B���4�P��zc�3�FRbݫB��1F�ݭ��,���G�a(d�{sG�\s���ߟ�e"�o�W1LX5[hm�-�n�&�#a��|��j+>fY�&�#R>��<�tg�%��i��IbN��bQ�����^��5S�^�O ����#�f �E�����r�u�-��>���cܜrvh:K� �֚��­��d��Yr
�(��� 1V�#2�h�4wy��CJʚ�doXhg2Ú�u�X��x��mi�C[� �Ɖ1��_����Q>9��O�#��z-SF:��Ō�I�d���#K4D���1#P��w�� ���X�6E�Q��4����<�C\��|ph�Y���?�^S�*# hš���D'l)�겨�+�B�mD7�Ok�{��T
���=��q��3����{a}9L�����+��Q;P�q�䷲��:bF�>���3A:�Op"V3�����_j���^
�}�>�*�{d!p�=�:�V�y���9����,�p.���Ʈzy����"�`|%�_�s23{f@$�/�<X�ڮV��Ŏmw��'~��S�������+K5�W¥����w�6�<��R�Ku��g�%,q5c�rv����B�9P'4��a��3�����G�C�hQo�:KTS�T���
(�tTB��w[���%�����Kod�����k\��v�Ϭ��W ��L�뾣9ea��1s�c�����*���&�������~������P~����i��B)K��T�т"{Y�$����E*��d�]B�%K��bH1c��s�>*w�<����~��o���}�s��z_��u���)��ZzH>݀b%�E�N#~f���/�öc�G���F8x��1=ۓ�U!ݕ�2��}zz����4w�[��c%� [��{��RsX��֣�����=��j�����qƢh �6���#��� t/���P�>�� %9�/���@jc[�A*�	Z?�lЌ$p���� ���3WvKK�C��}���k���&���MTM�ԍ�R�������c�	�M�M��g#�ؒr���/�������^�3��wk�p6� �\g�[}}S���,.O��L�]t���5-�������R,h�
��zL�lm�j��;��$k�{�����u�n��'�K�H�A���[ ���,큞�֫L`/�$�����B�0\X8~���,G��q<1"�Qv�))G�Ꭲ�֐�xGtm/�xㄢ���{<��
��^��X";����- t��"��M[%�"�(�l$@h�b�����^�&Z"|3&Z;U�pX��+>�0�q�=+���\��P��SÂ����݀�Y�
���.�m)a+I=\�!�9���t-3���y�}^�4�"A\zD̟T�6	�+�����$P�'�Ό֏[�n/R[���tfR0���~ ��]�S[��䄚��8]?r�c�R�v�ۅ4�f���H�y�SY)ܔJ�3���Z�߀���r��E�&�\
'����S�%)#��]�
>,�@����m���xuH�H��}b�)����[?3�NщGY�:*�>k�~������}	�&,�I�c��My���r�,2�U�zS�� �Ec�h���p���%�1�]��}�?*:H3@�"d%A:���8z8�`�9�.�5����j2�afD��-�}�s�ف���$��F32�3T.�d�/�lW� {.�gҙ�ek��L���|H{������SL)U��"��Wq�hv��>���ٽ`�u>�x�X3���	�+5҃���B�j�cMӯh->������3��=#ﲲ�3�Y^������I^g�-QO�9Z�F�Nb�H�P�|��h�j�� 0�oQ`��
++eԵ�$a�:����i�E�}�����ݬ�҇��^��+��|�����^b���󙨹B��ܮ���~��颤4�1��٪�8乣����g�pF�͌�{v�cq����>fQ���;p;�ڭF����UN2#+.��a��T�.:����P�#�Cm�[`�����b����0�����&�z�r��w���&uL�� ��xa���
w/P\�$��/���B0�9;"��<E�O��+񗀔�ϭ�]xxsToJPS(�3�Pw`�Ԟ�uM<+l�<@���P����-�4��fa����>b���)����9W�A��T��,�,�9����0;�-��-�;��J��}�j�/̸�+�xppP[4��o���	͝1�V�22d��A�0	�o>\�x�17�����fZ�qaO��<f����_��TlÂj5���|��]�ӣ�����UP�K����>��R�7���h	��C�� �A̐�!(���8��H��?�^���"r��՛��\V]�G<ʢƌ0�U�d��'���R���ۼwH�;rA�c�lA[���o�$@��B=�4�Q&��o�M�(&O
m5���xj�ӯ������hhh��Q�W�`t���m��
��^�G@�[ђ�}EVN��x��������O��oÙֲ�ΰ�W��c�Г�w��K�KY�V�[����uţ���H�ëޛ!�g�tg�i����Y
������m5���??�޹��;�D��5I�1�P���r���	��8��������Ef;m���AV����/�5Y���=���|Z�ޏ9T��N8J��JQ�WTF�Kd
�XLwml"N�RD�3y����Z	��aQǲ��8�E`U���h�^V�~F6.Di�������1e�_����jȵ,gЮ���ϫ�0;G��j[��O��Ǵ���9�������c�t�zVk�����G��h�)r.Q)y�Rla;uG	�uC���[�&��C/jd�k묃J�ރݣv�������g�OMM������d$�� ru����\��C"$��sEI���ݱ�djj:93AP�l2z��pt>Q�?7`��566f.��Γ�d��������yk e�.p�& ::�`H�ֿb�u�<P�nD+I������'|Lr4�R�"���z���7�����:�<�(���d�TjQvԻ�Pf���F&k*{F�:�?}�d��~�nv^^�q��\��J��z�E8��pk(3�n���U�ZC���:�#���/�]�����;�Eew����'?���0���$�)ȱ`I��p�ӻ�����e'eU���r�	�X�g�(9!ׅ�}N_� )�*3I�n��j��_62b9�r��ˋ�)� O2{q�Z	V��K6� �B�-N@B����;�����h�(����'͸v�IJ������Qjh��9�a���MV+�Z��=˱�;���	�F�x�f���S�^�����W�9��*E'���x�X��h�����e529��n"5�qP��yfu�q�h�(��y:�<B�ى"�������.s��d�קQn|b�""S��"#�
p#�LwzH �i�F[�Ϝ��b�A��t�`$09�N�-��-h��m'��Y3+e�^���[�P���ȁ��:���'��P*�2wr��5��Q�|^k��䖁k)F����ij|�cQ���A�ΊH�@��lx^sȷ����$���,9V6Z�9M����'��/[jǢ���h �g���
�20���.X4�O��Ԕ? ����~@4�(�`^nt;3Nq�ʕ+����4�l:�:����O��i#�:1��]]�2�K��h�_$��ODF�RM�ۦ�,�V yyy��Q8��.>b�B��{Q�>9yy<=��-�҃�z@J�WL~�*��(y�apw��tV%L�;:��]�e�>���Ɍlx�r�/>	�q.��nI�P��j�N�h�%����Z� �����OOO�< ��і{�m.qd|��<I��ξ�<\��zP��-�Z3�,�*ox�z�l�����`�qR%�A1�/��U���w�l�ێ�M����nL�wz!gl\BΣ�Թw���^��P���Įdq������ڮ��s��< �ffD"�z �̯��X��,'�C�*p���g�.l�P��J���:��52<�t���dN���}��8��|U�b��<#��lq��ÉR��uee]dQ�W�E�:�HTe�F7���������p�(;���m��31�|I��&�r-�)�?�&y�G�G[���ܪ��+�%:Rǃd��!��tE��|P6J ��;C݇�!u�VR-iH-�� �PNN���d�9��=��f�2 ��F��T���Pg>E����y�f�m� .�c�C' �Ǐ�24� ��fl)��vY��d���X~)h��Y��sή�a������|�}(>��{Q�i���?�g1��W��r>�"g���/ĉ��6B��F�x?�G��֝������d������#�p34�����2�]�9i��w�iy��pUj� B
z���0�;���I�*�L}\ 0GS�O �B�U�A5iư�I�+��W[��p�=n+Z`�t�%��t��2  ���ּ��"3�&�y����\��u+2@�܊�'Ze��t�9�94m�Α��<����W���UI~,l���l�~��&�r�
�PY���H)�bf_�͒N�n����{���ʪ����W����^*t#�Uy��-��.�� �g�+fi����-���]˕��F}J��'����Ӑ	 q����)3�]��w&o4I��U:� ���\W @f^ /]����s�,�s�g�L�A ��G��l�|G7?�B������=E-F�	W�Cu����%��>Q���'q�}�6��7
b���=��?커�|)��s�3u,��M
͐]�5R��. Zt����h���h��M$a.8/�G�[����֎Ӥ3��?��~���t�wm�ئ�� p�i��=�8���|/P�i-ƿ�o��|_�E[M|!��S���j�tՈ�������m�s�6���k�^|]�� ���$=N��:�ak�m�ŢM:C�k+���t��%d]x;��X�:i��f�yr�aHi4�;8 �'�ڕ �3n�l���j��:d[�%H�G�Aʍz�:u9�6�2 �[�읝�׃CB�"/��`|�"��o���7�'��H���!1n-z�����P�Z�?��M3���WIC&߃����-��\��V�M-�1} �@�%6�٢Fo��?Zh�0z�l��j$�����H@Z�q^`rQc�L�f"����C��w	�Dޑ�߈&np�����hk�;�Ѩ��?"�"��
T jcA���Y	Nu���B4�k�a�)�4e0;А$�n�m�ۤ3t(1sh��d�q��F�3���
��� /���{~���$I�h��O�d�����4��@.��@[���8�Id��O�r�6>�`�����H]m�B�|�I�=�C��t���y	�+�Ko?<�T�~�HBa��r��R6��d���}V�v&���m1��l���c������Ⱦ��7��_%�.��"�,�����,�m��>�E&K:�����NJ��Z��7�{L^=��,�IDkg?h` ,��m��rg���z'�����.�m�!����	ML6ڹ�ve�, >7�ٛ��Fb^���C.ߏv�o��n0�+߶��x��=�szL��k�zXo0��C����WǲnC�u4Ɨ���2oU�[<^�
k�G�@L
-��"�/������ )ࣻ�z�#f�v9V��ˋ}b���Jg/j�foG�)�;@O}���2Q�#M-;����o����t��ٰţ����^�p�����~�av�a7���׵�gU��z}c{8Z��Y{�
���?H럠((+�z�Z����X���R�Ro�M��l@�=��j���Hr���p�������t�Z���G���(N����͠�h���JЃzbY/4��{3���&�#J?�rX�x��=�)( �����h.�>p��5�}�d[�	�C�[�̀�.˶�`#�Px��Nxq὚�Zl��G��j�2|��4�FYqѤ�x�k���!��\w�(	��l����wD=Ȓl�KQ�QƩ�iF�tQ?�����B|�WZ��p�U����1G?�E?��� BZ'�pC�W���cA�H��w���+��*�U��Oj2��#H��Qf X̿ʥ
me�~:�k'ٽ6>����y���V�����c�n�`a�G�˒�BŐ'hC��=����ۏ�E�1��-@m=�/���y�=��_o��]�2t;�������7�:�ȫ��W]��&����&�����XLD;�\R��d;LQx޾�ǋJٽ�,,`ܾ�'B�>� JHȯ%�B�D�vy�Hn������]
�)!���*h�V���	%��9�`UZ*���� }�E��ހ�H�\V����Fk��B��Ae��-��p���<��P֜���-���`�b��<�a>
���R�IR��F�Od����&;��h�/�v�>ۿ�8��U���;3��p2�e@�9��+��C��ĵlXy��|����i�7�?���E8�e�R�)�:-2
���WU��d�A͜%� 3#�.�o��M6I�&,Id8PP����ޅ�l��m��,2 ��7>�k#�)2�3���\n����V�%��M"K�A�:G��?lʓE�ֶj �6L��!D�!X�j5K"?�ML��'*��!�����x�}(D�E��$��o6Y����ܩ�0�Qm�(�������6Y|!U,��i��Ń��s� ��g�d�	?����_�@G���^%�z L%�־>t��1�X"L�g&�5�#h�J��`�����mM"k������s@+�� �)|b���2�l��q�8(� ����o���J
Z����U��!��8 �2*�~�~�'�D9�k�l�P�O�L�l,EYYy>=���-Lv������.�る�N���2���h���[MF�j'4�����U���Q�ȫW�(D����%8Q/��;a:4 g��A\e��2X��!�P�l�������8	�ltm�0oy��}�B#gm�"5��u�g)D�R5zc9��fj�܃,�ލ���%g
X����{r���"�F&VS�P\��Y����,KVkn�q3�q�,3ճ��Q���#���`�$�M���I��#��(��Z��l�i^р�c�Sq�9���yR�@#;k��8ˏ0��j�8R�6����C'�)3r�t�	w�탩Q9�&t���A�3�P������D�X� 6��'˙7e�����ysy@�9몎GS&:���&��p}��l����_�trz�k����ʇ��Ҟ�e��������a�	�l�W �'eX-�v�AA��V��Ξ���g��x��V
�v[	�� � r��Q��Z�ʓ�A����V��u���U? �|N��0i�C�|��m_!�Ǐ�6��G�4Z������������b(.ŲQJw��%��?~��C���8��W�|$QN�������43434343434343434343434343434343�w�q���<u���lC�ֿ�~��FУ�5�ظ���?���������������������uf�~~MBn��ܯ����_��چ���������������������������������?������>�G���=^{o�^&~��f����=�^j��CU�_s����� �s����M0T*;)�k����e�{l�-����(f�?hE�����7�oh�о�}C�����7�oh�P���{)Nٖ�?44������K�]�����e��$��V..�*�84d�4MҞģ!���*>}j��M�������s)����5GG�Ԕ%Q\������;���3�ފ��U�Ј������m��

����_4ԧ�a�󶺮"�×����r����W-,�5�����D�DM���C���L]���ٛ`�����=��0�2?_�СC���g����KK���	+I��.�������!��Y*�����A���w
���|�l۩��.�MMM�?Usp�ɿ_��AMS��/o����������3�J&`,Ooݺ�05�[����ۉ::᙭&�c���>r��Jmm�_�P�����l�,���o����c-�Y)��_�4K��b�8n������\L�#Na���+�&&	��ZVk�KCK���C�n������ss��.,W�A�������D�\��l���s#����^�'8�')B���ו7o�񚿚;�[\W��Oo�k	Ď*))��:�Z�jK����oI�_}���6���J-Ou�BT�/X6�k���Y���ۜ�+�~-�ď^+Ak�K�� Y����`�~���F��ݯ����������!>�������e	?� �׺���v�������h{�?���s]u"DX�(���f3+N�#��p����݆�����D�ս;��� �?�����<����c�������������������f�uz<�����+^�Z��kU�O�9������������������@3I�N����hfhfhfhfhfhfhfhfhfhfhfhfhfhfhfhf�G����y�����6��k3R�j�0����gO]���$�����������������Ef��Y���lI����������������������������������a��K�͸����t3�<�Om��)�k���1z�<:_�����0���ן��_ZQ�C���~g~��q(����c��ۡ�o��#��[S>F'�w�Ȉ�����YgSڔ�&NR�g��x]�n�W�I^�������?VbK��k�8Y_��1�b߿<����\������I���&��C�ԯmR�>��'u����[�:�Cjgk�dR>�VM9��Yzʨ%�ӕt������`��<�K�/o0^��CJ%\�#L#����3n7	�N��s=�ǽ�=�$g���s�-����[M���0��8�`ۜ9��P�:��L���^����8F��K�}6Or���ϴ	��i�ׯ٧�n�$F��Ϋ��0ڋ��W���1�b��?wJ2�_ȴ�
���Au�i��j��ä53��P�ƛK�v�����NI��}b��eQs��.�ōu2jJ�bΓ	h�q¬]+/�f���_�t?�a�5�9V��n�����<��0ַM#��^k�����ޞslMY���γӗ�\=�Z=�\�?�.��Ql��7��3	pKx1�R|��5]�������/�lM.b�Q�:w�yg�x���;�c}q��2�[��#θml�����	��))���H_��V=���[0n������[���裣�>�^s�4X�Q��tgK���uCQ_}\gj�fܻ��fU���X����ɘ<+����>�"b��ģ�:^"����Zؖ/�tN?�4�)E]x�]"!|�Qa!/�+�����O�=���2*�.	��Y2�)H���fJ`�oL�bn�Oh}s�N���Wϙ�L	��å�"��7j9��v�:����|�c��:*�d��+޺�uBd0��H][b��㦞�m��������EO$�w�?*M��|׸&��{!ib�1{�"�R2��[(���J�n^���z�n�s���.3���<�)���+�����7r#ݕ���y%R��yB�<��7�L�f����r���0+���V���>�_I��z�w�i�j
��}׳˙V��#G���
��淙o};��,}&�^+��k��u�z-e�bo�͖	xx驨���aa�kn֕��A	����m�6��$�N�}!�髹�^���Fg�U������Wp��{G��i�ǟ�S�em�i���kv��ʔwŇD�ԾD�V^��-�R2k��1�|��5f||���}E�rf<ǅ�)�7��}Z������5�2Т�K�Z"�z$+e�1�	O&�gR�v��m��9�<��>�ֵ�	�-i`V`&��x�b��	�\��ӡ�٤�uI�K�^ζ3��j��S�	}�[R��|K��A������I��m3n~�@�1����Ƕ��
w�~�,����{V?x�����N���^�o��dۏGY��,u�fؚi-PîA��	V�)wO�	�:���#Ǵ��Vُ�7�ޙw~���ٓ.Ų|K�k�;��ҞE����7I��'?y��4��ŷk�s��,�:��'�u`��$w?�\e����$�`1J��n�bhӬ����)E��.V5f&�<V�e�����a��7j�Ǜ�$�l@RٓL��lϾ�Mn���Q����t5�z��c��������0`|��d�CO�I~�Z-�@�^�����K��|��S?���8i���`ɸ���c� �,�-�0W�ݰ�VD���ysO�7e~�Z)Z�|�˷���u�fdM��.ǙNZ\o�n��`��g�d�K��A+�#0	L�Wb"�`e5j��o��=-����������g���Qr!��	8K���c��3�{�D�~Tqk�
f���:�Im�I�Pa���'�=w3��8�E�k".'_?����bf�d��E����oo*�lN=H�b�n_�>��B@sd�݅I�	�%�Si����OB��'�|b�Aһ�仾�JT��SXR��1C��]�����H�a�_N���s���:f�;�Jr&��o]���K@d����g^�7��@p5x��h�q,�n��5>�6�XP&��7hR�0�b��#���
LW��;+�������%�`��.�`KOZj~�h�2��oL�x��(��ܶ�����!����Y�%���F!����Ԩ�hѱ؟a�az�8X1�[6j��{�2R����8so}��;g�h��}K�1E8�w�0;	O�>�ߡ+�Y���K�����Eٗ�kV�����)�0PcL��r��b<�j���k���:ģD��o�u����S��\��aʮ �."
���w��B�ͩ��L��|��;v,�^xf�Vgj��z6�'l�V�����J��F�x�V�MNUV��ڇoa�<ecK�,��y;@_I��L��LkC�TF�^| �ލ5\�!��,ӿ	�G�u�*��N�۝gGB��/�_>e.��|��u�����/I|u1핞B��~�DJOO�`�@)	�W������-+ȵ��̀�3 4����D���k���)%sۅ}����Lq?�ԩ"��R������U$�IO���gX�w�h��Y���yT���Mm����Cc��"	���3,t�RO�)�
�,(��W}'GzVa"#�G�U�~ ���xޤ��+�<�&0;?�[�/57�3��M������7`��2�S��v��׵�n�-X�����'���&b��~��Q�9��,[�٩~�ử-��zs��:>t����<���$KP΄���+<j�����J8V[���C�����o��>i�<�����[$"��C���c��8�"P{��*����o����z1�| L��j�a� aG;}��,%���[E�6��dq�����0n.T�~�n��P���uId�@ȍq��!�/��I7�11(˚s��� ԭ�g�\�Ԛ�j˨ߍ��5�O� NRϞÒ�>�)~�5���$�x�n-[U�]sGv P%�ؙ�w����`)�Գj|�9�pP��ɪ���I���^9ܷ�| Z��X"v�
���w�,{O~�eq՟_�Pg��D�B��Y%.@�|gd���@ ��~�Fg��n?����r-O���[��Yt�ٵ�Z����S�e�޾#�R����� ]5��X�2G.�����Y&�^,��2}�!,.�ڇ{C~U8v�TmH����Kh��:��赶ɖ�`,<�9�gLG����ٟ����r�	�;s`^~_�(%ٓ�y޵/�Op�A��#�}nLkN��=N�
�yEMz!��j���[�u���0q\���C8N�ᩑ6Gbe��;ؗ��k�8�3�6W�
0y��o��ފD[����._M}�<�  F6�_�4�<���>��u������K�/e��d�L&w�9���&�����o���M 3�7����}*y���R9��W�K�rAH!Y�}ɡ��έ�v�<a�Ì�ɣ�B6�قxۀ� Ap��K�Ew]g��H�9�y0���ܹ⺦(n ���5����&1c�u�+i�;�IwX
A�Z��dM�X��\�8�kv����7x,���D±�OAL��k���8R�Ϧ��ɛ�~�q8��'Y��Q��1��)N�q�բ+>�yӏ{/�F8�#�a�!����%�ևv�(�L]��Jo?�r̴M>�������������Y�c�F�%U��Ȗ1��@ �z� �+�Kl;�	D��ϔ�b�*_ש�AMǁTn�lιw:���?�|�X�t�'�_��Q�� �S�/��e���7��A�Od%�0�����k��Si�s�Us��Jl�쾝�S�6�(��9�J%HY	P� J(��P�@L�V7����j���[��mG�'� ��s�y����_7��a�E����Q���ѱU�v�}��!��.d~�����_�
1�ߜg{����xϙd�g��B����M��9�Ŕ�i���]kZ[L�OL��h�ť"KM�k<�uw T�W#�Q�^��z0�GJ�i�?n5'�Js���d�DZz����!��0;	�zBl���%�PE,@�EN��+��շ�Cl�����1o��)�OoS#�D�	ؖ�켝%^^�Δ�t��Q)�NLt�������<�.�]Wa\�ԥ�U���y� z�xw��V/ѩ��)
7��< /�휥�@�^O�v0X��ph{	v��t������`�BM2��1��
EV��D���c^�߷𙊦�
���BSC�a�vz���|�э���64e?�
�]�t�<yc�yi��8 $6���U	LqG�XN7^�$ۓ������F`�k��uz��2W�N��n�����z7�x�� ��J����I5Q�|X&�H��m��Xǰ�>R�X����\} p��ݷ�[��B.䰈k�秓F����hyB0l�����.�\�v1�z� ��21`�	3�r��O$�A�(p;��| ��v����|����i[6����u'k���z��6��= `$�MZ�L�	�tcfD�-�/$׶�?�ͪVf�p�����ƈ��7��u�6&�0h�nI6mĵ��F�׃�<GI�Q��8֙㨌�<<54!�E]��QJ2��f��r���`"�|ri/o�-������0�Ï�?Շ �U�� �tbȾ'h{z��y�׵�O��5�!�+/��ײ_ѫ�(�涛���X�wgt���
�lV��̫�)���ļ`�ٲ��sI��}07�ȶu]�m:�O�ɗ�?����|�/v�B�-+�m5~<R�+:&�_W�?�����P����C�Mo��(%5�S�@��^��D��zsu|MD�5O�R�`f��~�N}�qڈ����Hi_u�\�C�������8���~01���,S�nɏɧ�-�	���f񖩮5"0`|�d���G;�N_f�-�I�h������[.��<�,�g��.�s�?>�19M�Ʀ`" ���|�wK��%fU��{��{��j�##j�1���y2�Q.�3lL� bU6����Nu�h��#��/�x\)�j�]���pג��R�_j�C��<IN��xUK����9��œ�J�"#4/㊾�tYe�ȥ�L���Z�0m���*V��W�]�=��M�ZR<Yqk��1=��4vz{�?D�D�];r�[x5�l���Y�\��gno�5@��l��!up9�#�u���5ҿ��*)��=��3j�[m��yRZݶպ��3Ҡ��~���3w����!=�e����/ =�2E<����݂�@#c}.��;y��A������)�9����)��)�����Q��'g���N0��+0�d������aD����D���3�U��B���!�)7*�>1����<O�'�|����RZ��R}�]��9i:wcW�W�@�n�������y�"��T��\����ǔ*� ���Ə,a� Z6h�ME���!�<ŗ���� ��Ɍ��,��\7~�eV������� ^Dd�9�d�2� ��uGS���7I씂�yѶ�ɺ�ꆍ���F�0���oI7�z2�6��܃��c�،�����JtS	�3�a@Z�����<?.ep��"P�H�3��J�ad��G����z��7/P$1�s{���C���u)A����7l�n��ȴ*-�b��2Q�|S���WP�����}����!��Z������fE1\�c�Q�s3޲e�ʯ�]�׮�Q�ӯ��|����yo���r��	���)�b]��(��ȩ��t����D?����k=���'���C%�6��T)�s& l�ݴj��|Bj�@��C:N���l)n����j1�4�:Q�U��A����~K���RM�0B�6>�jW�ɟ�N��ߜjHc��1�|"P�)�Y>w�z#�5��>��㫰��/Dm h�I�U:�nk�4�RغR?�"��j�z���U"Ĉ��'��xs��n�fZ��8z��<����֖����7��.-�u���;�>J�\���6?_�\*W$$�}�M,LP��>�����r��@�)$(���Iw�w�j���vW��,Y�<R�A��<7;c��S�<k� ���h�o����Yny�i򐪙���D���7���6�%�����ٗp���9O�f1���l)�z��L !�~b�*ي=ɳ���1��]��ż���c�	 `a����%J��5�������r�a�ωZyꆰm���r��*}�pWy
�6@݌z���)ڀ�C�ɩ�{L-�GҀ�6Åʧ�A�T!`}�#�zh*���OJ���!<�K�6��0��?>as-Pj��q�Z�:�Z�b��0[���_]�,��iϿ����^>���ܤxՔ,lƁ#I^N܀s���A��V�=�>�6���;?_�����f�T Q��w]{��L쭍^��=�1ثUw�k�9�����+��&�R_W�cB��X"��Y�;U�ԝ��Y��"-��S�p�6� ����l�\��x�S��� D7$��pe�������hD~����b��;���7�������w@f��{��L����d��ҧ�����{�-}3;�WX)�y4d��.<�#��H�s~�x�@��-��3'"%�Č�t}-OΎ� ܷ��`w���r�YM^��<��j\=��x_�I�y�N��R$��z!�����jF&:f�p�gz�OP�^C��P�W����=g��x�<c�����W��Ӛ�aq/"1��}��D� ��o,a{vP�*��B@�|�s��&[���C���s�a�Z���	-��^�S{�@k��R�m�K���Xc竸����O�8�ԙV�A �d?�*FJ��I�F� ������b��U�4��"Q"��	���a/����tL����C.� ��۶��%�R�C�QIԄ���!H���o�����a)��Ѽ#���S�as�ar?S�D�����3]�<-��5�x�x�� �3�{4`�_Xy&D�.��m�1 �w�Zt1r�,�L�ާ�9�����څ���P��)ӱ���y29�o���se�IC���c\S_!��{
��{������nkQZZ�,MX�É�T�9��.?�Y+�5~+r�9���0��?=G����1I�������**�Qؼ��^��������'ɢ�,�,T�땢e=�r���wu���"O��`�I�W���>Ϙb�̏�ᝀ�?�x|�\�h��a%L���Ek�v�D�_[�0;r7$j�<�Il�1���H_M�0�#�_����u����m�R
=�����U����[��A	{^��:��eP�J½DT`�M�p�rX޶nD�<��芌Ɯ�{LɔP��M?�c������m"�6�p�V��u�O��H����P)<c7�wm���Y��W9�κH�L5ɛ'�}z�P��������Tt~�[��\�Uta�2��Ы�����_���HW�żm��3/0J9<w#|�s�(����V�E�??.e)	ң���KU����/���Mի/ۧx��;�g�˜V6���,�°����_O[O8~{��D�����^���v��ʌ:�Yrg����~�.n���?���n����>����v~�ڣbp�u3��Y/f�X%���A:����<7"?�'!k0�5piF�����@d���v���w&5��l~~�z`����9`E��c0a:��5�2/��X���||p�V�?%Ձ$V�h�tWZ�	:�Z������j/%��ջV�JQ�����Ό�F�dl8"���Q�{�nES�E`���T�_ݠd��H�є��ip���x�*c�k�L'������d"�%�^^d ��%2~i<T���O��gA>�;�[��WD�}�x�
��Y�kd��������b�Xr����CW$��3z �L'��Й��T�)o��y���4Xl1��a.������Lԏbț��]��9�uiOnSY�P��dL1�?��͙�&2M��$=l���J9���՜����g
��^g�Twi�=�j���m>;�#	 �@���g�@hJh8 0��E)�i�)�>�\�D�*֮x�����}���OB��ve?�#e2Y��ԗ[uK�U0�$@���d�a��b:��+���//kx���L�瀓�7xN�WK}��j尻1uA�=pc�[L�gY|7��)o��_\%?�п����J힙 �$�N\L����~x�2�p�u��� ����s���]�#�_��qԺ����\�j&�]��~K�tΙ�'��
�F�F�OD�Y��'2�e����j���]�m�޲6q�6ɆLSGۆ�U!!�z�uS'�{�ˡn�nɛ����!��,�_c3e^��|+]G�`0Pi���J(k���ᒒ��2��tU���qD��Zת3 ��k~��Y���O�'7O���3�VH�#�X�����I��wQ;�L�������Z�z�9�:�wo�Y��\x/�a�<����5�֋G#��U1Hv��^"��{=F����y��7�L`�X�j��2 �����%�6Q �Y�Zo	���������q<�pߕ�O��&er0��HM�`�2}��}��}�=5N�ZF���q/��$3A����:��NU�+of�4���3��Fe��0C�6DUn�g>��6�<L�	�F�US��~��	R{��s��]G�+i� -)	�����=��>�r�.r����b��mg�6zD�t+�V�"{�@/��_�:#Q,�*PUa��Rj��]�y� z@�c��AN�u����u�޵��5����h�}�+�t��e
�	xG��6(y��`����Bm)b�K8Vk�,C,]�s����Q��H����
��,���.Cw�W���M��8N�у���e�̙h��z�cn���m�Q�2?��|k��g�����|��P�yX��=s�Jx��n���v1�@h�h�|ћ��Y���z�����R9���	�B��-�N^+�K��c��W�ok��5f���o��˩1	��+k�}u���`���w�>SP���@l��y5;C�L�Qi��Ә��������ڧ������p�et�
�%��C
4;��)B5��a�r���^J�GW�
�|��'N���|���}�@��7Pz=���S�#*HG��0B��j%�ڈF��j���|l������/��+1.�7��j�}%O��t���zw�S8�����o��iݿĉ��-�x��.f�=&�d�)�c�]�'y4D��p�S/�������Ƈ�@P�[䦧�$���k���e�B^"��t���������7�#�1�0�pL�M*�>	�����0�(��"���ɞ��F`C$S ����p���zQ9oޮ�� '���%�9q�Jҋj|�]�N�Q��,(Y5�#�������s�x���lvj/F��ίK��	֓��?Jb�:��y0at�Gw�9u�NIn�)1�Q�}���=�8A.Ή�g6>�*�]U�����d����]*kXo�諏S�WkI7�R|cҚ�n䓐$�u҉���s��V"~�u�)!��ڗ3\v�|nf�Ӗ�O���g�b4�%w1@%y�o���0P��x�&��G�KU�E���+�1�"MD��U� uZ�غ�f��Oe�[Wa6~l�ҙ�.�D@�?���sq��	@^�[aJ^��_V�\iS]ۘ`̉{j��5:��v�#ѹa[`]E����!��TQ�y�d�ʧa��I%� <�a�7��͵�`#?ηMR ���c;�$�wE���%�m/*�~���S�T�s�j?#�;���=wԲ�B��٧�K��2`�r�Cz����|�K^`���c@�ɭ�a*��X�L~�t��EC��u���ɏ��E�)��I����)�Á�t��sģYH#hnL�0����#^l"P�&�]�N��)�`Ψ8�+I�o�XWv��x��Z��-G�Qെ!�U�U*�����~��&��)��L��7��@H_n�;�[L�ݝ�إ�~^��	��:��*����`�GDN[�tM�S�;o�P<ִ��� �>qi������iQ@���p�c��d�fW8����'�2<������v.��
�^��x���P*������cM\2Y���k���Ӑ�	���g\�A�x�RȈ��9��X����,	ԙ�=P��:�R��<��	��:�ï��ĭ���mZ�/I���.���GB�������]�g��̰��m��&��d����u�COA�Q�r�PML�铤S"�Y�ag;Ry�2�/�ݦRJr[���� °"�8��p=��ˋ�4�H��rԗ��>װ�[�pz"������إ�S�n1��8w��=UNKM�PF�&��ɀ�u+���?��.Y��Wܩ�1q�ht�J�}���L��	�:�x�Ta��9
ArOD�C��N���d�Z��3�y��Y/��Ρ�/��Ô)5��^N}�p��N1ev�������y��JK&��5{�1�u��o��<��}�������2�9��m	Y�TL23MV�&��6�q�4��y���ֽG��]�v�7��%�?�)�ŗ��Lq#�ƛ�-�c���Gs��Z�l} �7'�L0߼�:� ��l{�џMG�s��DUA֎Ut�-=z��s�Zc��;0�T �~ߟ+�2m�m�� �)��`Oܭ���l��ۛ
|����c}7�; �R������ɴ�)�8����}��W�Y�p��b�Ν�!f��S�R��I֯�zjP�,<�4��s�õ���0f�������͝��"1�[�!<��y�g�vU"�ДZ?�	��ij��B�M� ���<�	i��Ҍ��6�v�����̖\���`��ЁdU�8~V?�8��/�����Ɗoc��B̥���;��o�[Y��0c�����*g�*s ��7����;��a��GO���r���q��ۧ�|��pG��
a�C|lu+���",amY�ȸ�MZ���V)�ó�����K�S0*����\p��`~<��vT��0�x��`FOr]S�^Z�j��.<��dB�o�����@���Cޛ7]���yn��2��À������X��'dkRJ(oN5t�s����(���I��ȘPݮ������+���4�ѯ$v���͡���K����l��w %�� �uP�}�(���QPV��r{����lF���Å�|���߹��94���\'��T�����������4pGo\�#�@�	��2o�Ӌo���%��\%<r�yq��|#�tB������`A�{���� ׮���T���f4���,��Ua�U�1)�gH��F5x�n�@l0��C�����lB�T<h�\�y??\�p�x�K�`�7bS�_=lj!XV��:O�~��adU���@�x�b���4y艴�}�7��v%W�&B?�Q�-�^>r�� ��
6ė�V��c�(ݶ�i��> �_k�J<��$�� R��Ov���5�睙Vzg� ���4@6V��Evm��΍+)�����ʰ*��}0TE%lAJD�AD�F��:��4����4H��Q��HH��C��:μ���{?��������y�^q���uo.� L�?�޶LZ����B{V���y�Z���A"�>ZV�^���Z�� 꺭��=�>���'r�=�������e�����\B��nS���N=wF��6��J\WW�;�GӟǠ��r�X}<�����aY�6Wҝ�%f�Җh~2E�D����|,�݂�PB�$F��!mo)x����Y����~��Ud{bh���Ai��m���<)h��x�Z���U5"W�d�山�̴$�2���aW�Q�����Q)%yk���L�dG���9������X)*�e?�$��&�[M���vH�XZk�����;/�0�&a�Ԇ�-�6�'I�F����D�Uu�T!}T7+ٰ!����H��^m
�����݈U������M�=��}���W(`h�]�O<E4{�Q}���|E�65���f�����	8�}S�j��>Oݟ�����Ǒ{9H�)_UUU�2wJ�t �B�K��N��T;��ЋQX@�vJ�"��[ﺩ�p��xzG�����Q����v��sKr��$Q>>χ��/Z�ν����s�?]���>������[��[c���(X;�����j@pp�rW`z�X�P���u�@���7N�ũ�ӷ[G���\؆�K~��!�.��h�9��'`�`��ro��V�����>���+X�ئ����q'��t�i(U �d���l��d�*=�r2P<����=����㸽���9oQL�@���~����df2��(�&�o�\����}*^L3^[������Ÿ2袲�ߊ��f�f���д������'<yB��g*ܡ�K��_ƺ"E�Q(W���c�ޜ�d��m���8�S�bq��p�P����~T
 ���k�ԫ�?+y�������Ȏ�U���')�'��޷��e9������dd>�����Ɛct�ry��;�󓝡��Mӏȟk#|����t�6�ndhe��=����G��+C��-�(�颚�d6*,�=o����˝���k_���K~;��
��u�Ňm�,���i�`�:y�:���i3V�����G�?�D�@:9��w<�ۗ��7�/���WR�`�G�9Z�rT�!�E�R���!;�Xb4�Q݀2� ���F\�D�<����kǃ�tTX����oe,�	��z`oǳ��E�9�&�m��%��n�n�N�#LQ��u$�~�l�Ա�;��:mJ���p=g:o5Yk/�Ll�m�y���5}٭�$.b͟������/J����8�lN��X���|�/��n&��y�	��S�{� �x�9��˥�8'���RQQᇉ}�ݠ?ޖV�%���͔�l�-
;�����i�
�v���bn������p����E��`O9w$)%�a���%�j����@�4��6`�U$���y�IBQ�����2����"L�-�P�Ț\��ܣ�(�V�[�1�����崺�ls:�(�_�X�.��ȸmX��8N�,^/��	a
A�#Q������}��CT&z�3D����>J��Ӹ4�O��O�ޘZ��3�n��8[n`����C����,MZ4��hks��(n�`˩q�E.�gt���O�q�] {�o���u!��|���G��(����Gx���a��|8�Bڝt�dkyK�T�M%����3�@{�]ۻlw>����1�f��ma�,R"���ʃm���
@��1Xa|���Q���-}T�{��+iU�0��Ǩt�"�?���2�!1��ȳԯA�+���n�#�-��E
Ԥ��jQhSRR���ց���#�����+��+X���R� ���C�3��#���4J�tS�^�K��䫌��E��iW.�&:iǾ�[Uc:��olh��QJ���iݪ��zw
uzYq���Ha��O$�T�M�^���Z�3���ݴ����2��_����%Nq��Ȣ\��D�Kq�����}�R�-!�م��1���qY�� �A淓pq>�.��U�{�m-'��y���-�x8�6,J�B��$,�ݶ�A���mrѩ\����5J��8��-4J�c S�Bq��`�	��A������"*��W���+X��ϺI�,@GDk�ಔ�n�B�l�3����#﮷��[�&�A8I�;rX�Խ![�)���2��6�'��FG��&���Й�3������.�V�tJ�6�k��_5ɒU����y9�kr)�t)_���*������')<�rk�A][[{WiBJ\ܳ{����j5�����r�P�m����Has�l�#Y���Y���������[�}~�>
��){q`���.3s5o�/&��\?T�~-u�3��=�ٹ�����V��1E4�g~.Dh����νlnw>��%iX�����]�P���Vqm֌���� :�P-������MjP�n�� �zW����+i�
�:��,J�ԑ�c�	r߱p��"DUۉ�������6�m�p�8Mt�z�ʤCϚ�\0���Fo��"T���#���m� ���n�d��l����s��%�)�ҝ.��'�,*fAR�ø�j��K�aK�VI�z�Q2:������ ptQ^*�k�����N���gE�I�or�ռDx��܎>��r�1��,H����&�Y�a�C�he~�v�ඈ�G,��<��o=�sڙ����(��79,C 3/BYD�k��6`9|�w��!1T�؄~�g�<�A�h7��G��IC�E��vjt��C���*��6�i�]�_�"t� �"ɯ�Ґ�_Od�x��3��1�����;��ӽ���Ss�#��,�� ��C���+W5Y�α�&���{��I�J&�wVe�j��*�}���p$��'�l��5�.���J=�@	�*�z�u�.�T��)����q�G[mv��gq�{5��	u��01kkkR��<ڴ�\��E�&U��2�kӐSb�n�5�)v�D���_��D���3+T/p�e,d��r}ց*������L����ߢ$S�7��D���9��G���8d�H���#�'V�b	##p�`$5\N\���J|���K�}3o���2R�I:�P�{��:l0�"*<�Q]�{`�_��UN�y�{p�)��ˈ{&lI�Ǘ$gd@�M~�3W�6�,H��%]��Qp$���l���ܙ|��.������(9��;�����E{����2�����#(.�xP_4oT�Yt��RR������G�T�ֻ�����;����83Q| �Z�=�H�؈��fp�NCdxܐ�W;�d�e��4m��S���Dky{4]�ۆ ���B�t}s���w��k�9��%	~sZ����Q�埶���G�=��P����EЋ���
�9jU`
�X����dP���q�4l�w�hB���B�]���y�S�:8�@b$�Xiзi��#ҫ�R�dyO��B�MhSaȼ�,���Z��(���R"�|(��g���rT����
�L������D�%y�M�.!|X�Kۚݔ�i�n-v���?�B�
�H�<�Q�io.<�y'L���c�QM�����1�8,h�j�����U7�)�p��_� j�}4l/�d[��6����፻w��?p�~�(�7���W�&{��3P�a�H�N�H��!F�V#�}*Vy�&z��*�n����	���.4��E������B}ݸ+���0�18�k�����-��'_{Rձɹ��K�9�}'�	2Șc�S]yd�r'?v������������xs}���$v��������H����/J1���NH���9��#���۬Euyv�C���	Uۄ�aQ�B����7��u�$��`ƀ��|7�c��.�o��}u%ݩ��9�7��Q�͓,��ģ����~i��������&� �}e���nk5c��
2�[�y�q�'�J�цnƑ/L,$��,���	���r{Ij����.h��j���ЯM�p���kW�],�U���Z���!����:��[atRӿ�	Rղ{�V�$q����lG�����e��K،r֌�C=[�˘�޷4\V\���ʾ��2��Y��m�O�C��^Q�eOT�=9��p����wh')�(Ǖl.控���j{IB��7l|my�ע��� �c,yuO��02�u���u�ӅD��4q���g�|�N�+[5��ų�	�r�=Ga�)�m
�/ާ���.�am������TӴ�=��H���G�c��g{5�ǔ̸qR�1+^�{{���|��4�s�i�]F�
1�����[�=[�Sn�y�C��4�ɛJ�u �o��8b�(I�*�[_��,��'(�MHA�����0V���h67��D�X��p׳���;s�e��*�h����*V����v4i��[��ܒ�<��Q�d����K��*^��$�$tP���F�Z��?�w!�|����Q��P�c�ko�q���ڌ�^4%����$;U��j[���)���n3�򭛊 W�G�$�w�q��f�OC�-��欯g��C:���4�-1!��+�E����suat�ڕ`�X2if�ѵ�	}��Ӆ��sդ�,n����֯��X[��{�����^I���_�t��u]�*4:\�uE/�v(�r��v>� ��+{�L�O��8M6��i�d$��f4R�u�S�'o�=[,E���|�	���R�f�ȧ}[5_�W#�n��@�j�" 8�*��ľo�J��S��g5��P���N���s�l�/I��A���(���U��{ನ�r�č��Ǐwqu�oއ����[}���Ћ���*E9R>P��a�g�`�S���B�5x�w/���xs��$�W�o�Xב����v���
*� Й�s�'�7�V$���
�~��6@1�'����Z�*�^�r�
@ml��B����Y���j��p@e~�H@|+����jј�2Q��X
DKR���/���o�w�nd�e�>��Z��Az�����W�л~WFa��t�䂛�zCp%Ɵ.zn�γ�N~�����
�\�We���%�� �j��9���е��ܙc��ő?�����Q�N��t��;Z",gpX�&�t�z�78KP��_i4�T��$F&BJ�jʏl}��d������R�b�Q�ɛ(��W�� ���������9���(�x���W�$�)��+�a��z|��ݎ�C6���j�����Xe���~��UrC�9P��pV>4O����1r_l�Q�a��������J��k���T�x:1I���h�������m*�����h���\�ߖ�+�9
�8�~����U������dr2R	9���<-���~���cI	ۍ�8'���0XD�{ˢ�E1�O蠢�I�[mz�#�P�ˊ�s���/�Mͮ�RFY��BU����F����Q�x�J�gOz`:��12�J/y�l2fv�R(4����+,S��qY�u�%����X��a��k.]Fh�)))�_U̧�м���Z$������9Z�(����4iw���E���-2���kSNmۨ������W�����z�p�˗/}Iu���E�k��	��x �p���զG8��<��
�/-����*�����ĸ^��3�:�0�s3Qh��S[x���	�R�V^G���z��������,M���{`��?��AV,��4��$�ƒ�����`�̄`6n��o
)M�kS�J�%/m&�KLQA����݆�6�b����V�ȝ�_|C�D2�E�ݥ�;��ew�vr~��m}����u�Kp��I�(�W��~{W�q'��D<vU=]�`��p�AN����T'��i`"�B��%���	�&�5w$*��\�?����*����|�������0�GƊ'_A���J��m�?$?!��q�|� (���^�'yA��\�Uy�ߊ�U�]�,�-Iz
���p(��� m�0?�/�"�E�o&��v����R��M.��8��c
*'"�w����:N+A6\g��K&
ORz����ɮbߡ����AN~O�ڠrN�`��w'�#*]��@��͚0~n`S�l�z���&G�岁ő�h$_��0�
zU�WG_��C��.T����%�Dh����EZ+H,We��Zh�/�k|�ȇg[�J7^]~�B�R!�f�	�[��_�x���vLD%	f�4H��� �-w,9�Õ�uӗ��s��8��L�����d�H�=@�6����B����n��Q����(N��p��=�E$�����Ч�*���!����R�v����%� 0�,0���N<tmʪ�͋3�V�)S��CE_�����������<K�K��j*�����}v:��k
![��$|�D0�u^/�$E"��lSpeJ$]t�&�]��p�׿:�3��� p~J?fکBks��o='�gq0�µ��_�)]���ʡ*)��Dʭ���N��dҞ�����Q�$�ģP�-�x}�S��f�#�n���m��g$zU�0/%��.�w���G�QTC��s���LH�'��c�P.u�(���Ow)v@}�����/Ov�҇�Nu��kk0&%5�?J�5��)�ۤ�J�wr����}����(���]��}f`�<5yp[3�7�(�x�aw�]9�|ڍ"P�
��7�S��D��@&��k�'�ޫg/��g�0E`�}�`�1'�[�"� @_{���~�>��BسH�4j�ҽ	�
0��	G�";�YEU������������.������xA���ܓ�����3����Of=�f���E���f��7���6��'SV�#_�"|�
�.��a���՟������f�L�j��!Z�Z &�F���?*~��Y����7 ����ZYe�r�v��nKB�4��F^ǁ0�Yz76T�?u���%Ú������k�/��u�]��%_����6��F����?}1������W��I}.)�w����I�p��,����vscD��T���濢TN�*�����L�fp�ޒO�����n��I�»�_�C�w]��j��$|B ��I����}5��wX�1CvP�t�4+�RڙP����iV�}�\�q#�YA�z�6�&��У�nM�4w�\�A�"=����`l�MZ����	���b5�>��i�i�x�l�;`:�\)���,�҄��̭С)�_$�C0S&�~,����;�� xE#�h���%��g�͸9Z�](�3���%�F�2wJ�P���Q������w�?���C��hC(t���-���W>/���e/p_`�mP��xb�9�����kmq�g'�\˔UUi��L�,w�T��ڽ�L�$��Z��GX������|=���װ�W~�t�	'�53�K��OǇ���@>¶`�HO���l�N8���~燠�q��Fy+�q�>]�^l�. u���1]#6r�Sm���]�ĵ1"�?q �H P=!�9?b�84s;I���$�<��`�84N��Ipf�o�i�Vf���C{{�Yh��/EH:H3�-
Jb�3 ���i�]���y� ,��ԉNK�����fR:-]���I܇����o˼��fz�8|���k�ғ�ߡ�����w������E�������1�>/mn".�b��M���[o���$�M��H�XU�}V�%�D��+z�O�xcuQm��-A���@��v�C7x$�9%^K^2�.v��=Q.RĜHy
(e���4�3����M "Ɋk����Z,�-���ɷ�΢T��"����U�LY�Q��,=�yE7�����J{�$�Z�����z�`���$��SG����"��<��o�jO�1 �'�_��<��Ff��S2��	�L|�[���X3�cP�4�pp
�K�K*_W�߫�8,�}Z��i��B^�fj0����'�}}[ST�2]q$�@+:Pf��q�la�^�@��$�eu�v�Y�.�N�O��u��Ձ��Ib�OfX���~��;��I#�o��h�^A�U ��;~<�%��\Gh�.��ʔ�_���(�t/[����"�oM}���'3��ևIA�{���Q�7�J��(������:P��ȌC/�Y�.Xf�-Mm,�����l���^�����a5P �*�-�G���̎��ߘv��ZB�-��C�-��;$���V����H���?�r�xڧQa����va;��⣉�Ʋ�9��)��I�Z⼡3���/"$`�E�d;���9��i�Gi�/��F�ʛ��I/�� ��ؙU��Ѳ?����<�K-c�x8Ҟ��ݺ�ekp�r(�~�D���|Ǣ,��P�$L�E��Q�n�b�N�Vp�p���������L��_�� d3y,H��X�_����IG�wEQ����~[�~hY��_�� ����Ȩ��<Ro[�䗭4�.�|.l������G�nг��]tf$�33�dW�Z��i	J|k��-"Sg�+�h���R�O�M-[���\.��"F��T�� ��؉ăo%��aB��}��D��� <^=�ec �BP�?�����04�3ͦ�N��㿖��%4e��b{�Pq	�O_r��K|u�S.��wlX�U��dM�SPL�!�G�Lګ
�Q(�>�'���������t�W���i�A�H[��Q�H����<����,�SӛF?A���`+���d����O�C���?hp��@�E��������+�C���+�����~�}�Ԍg�Eޣ�Z�!�[�A��=�@+�!�']��s�f�IOԊi#��j���0��L�GK�,'�N-B'���*_ PTP轏��FlWή�˭�@j�&���K�!�,¼���(&��-2�&R�h>:��N&��V���V���`<3os��|�^�Am��m���y<�7���n	�"% W���j� ��Z��jn>$v�����B�h�c��k����r^402�P_ȫw���V�7-��Nu�����TTcݛ몹���'�r��M���_��ZE�w��8nV�&N����]<	G�1��l4�h���w��P�M�~}���� IR��
_&&��k���$���N��e,J���V�S?�g�
��j`�����},����˼h�ca�l�+&ʚ(�S�é��pA[������� �����|�Ē��L���K��ay*Q%��n�I�2�d��O��r��;Mv`=�e$&,���S�>�o��0ⶏvx/#r ����&g�-�CmM��#��1=�5d<�
m�,j��u�X����Da`�f�\;����wV�/w[����Ɩ��q�����p���;�Eq@�,�c5�$"��@v�Sߞ8���e�~m�/!z6d{T��ŋ=b��ޒ!}	�V?�0?��[�l��W���Վ������ ȎG�j�m�����u��ڞ�[ k$��<���G{�F,1�֡x*��7��rP�ٲO=ȫEN�D
�a��wܾ�_�=�=.HK}W[�r������=i9)���,�Fc�<HN�,�T}�M�|��.8"1�G��.[�x�3j�m�<ݝ�����vh��.c�3�$�!Xz
G�pv]�k~ �00=~�r+�2K���9�a�Qbg�?
T�(��Ƈf�v9؂^���o5p@i�������?�hG�V(��/..�&,(��"���tѭ�2�%�J@�E}��q�wW�*T؁7��L>���V��Kd�mi���$���uP���:8�]�/dAo�#ha\�J�e�-Dt���h,O�:[Vɤ)�����Y�(�-��P{Gb� 8�k��w(�^�- 	^9O�[@T�o�p>�UFĉ�#@B��GP��)�fr?���F��M�]��S����$2$�����ӸFc�\���H�tC|x��ʉ�S3�G3n��>D�g{)��m�����2�ƔM�SR�os3t����L�"�Hv�q�e�Fd�EIm<8ӧ˙�e��Y�z��@��Ȑ�Q�wD�����������|��ի�����xM5s ����{���`n}ُ'� ��y�]#^�q	E=kE k�:�K��A�؍���UeB1�'��݉}w:h�y�*�7p���)Z&Z��Tv�>�&rQ�|��씮��m!�(�;	I7y���'J�@��n|�w/�~��fd�����}Q��r�MÌ�Q��M1Y�9��-/%S�˝�P2/X����J5����:��0��{6���@���e���P��Lv����Ǥ���1����5>��MP����/��-��;��ul�����[�� �m�����'3�=�P>����}�\�zc���|��v)D/�)��:m#��o�t"!57x ����J��.s�]�h�vW�����8-��Q�)�n[�l��X.��S�ٞ�I;J��O#��Rd��*�n�àqTG,�0��"k+ig�n�;����.�~��x	��y�wrΔ1�!������P"���B���6���mG_=�k���u��}�?]���.A�����P�����\��lT��N����І$�����J��o]}�'���ƈ� JeN��Dl�E��D��$ʞ����NsO�q�����s����R�w�B�`�d��@	���\.�ڀ9�F��J�㪻�0�@�=�i!�iY�S�4��$(tW9PʃU<���8[�8�J3C���X}�|�`�%����ȕ�EW}�a.$�Gδ�/��;A<Rx����+��,J�蓩�!�c��# ��cQ��#�\�޲�Km,Ε�CI�^ȦЖ�;�Z�0�]���H.<�b�<�lz�H�gт����(�5�P��"\T���w¬����Z��gc�gs�ײ[�T?k�J�����uuua���EA���{� \����c��o���z*�e�U@e�f����mF�΂@W%*����6��F��@B����_�@I�Lu��}��mɧ����K�S�_
�6�H�?��)v��T ]�9p�E�w�Yì�q��
������,`�A���OzE��?`�΢�[�0�\�1re��֣/��kH㲷��[�&�vL����J"��� `��~ًr"�`�a�T�O�@2ǣ;�Ӊ����$�p+�c��U�yC��g�"G��E5�!..N����Z��� ͂����G�GTAQ��^+������ظFQ�L8Զ�c�3M������u�j�G<�1�kȵ�Qm�;,���Drᕝ��c;��-��3�!�L��J��P� �����|$�~�u<�hA�s-��q��~����=ƾ������H�p�B�i�+�r%29U�����+������.�Z��p�Cp�U�G���-�_�y�=�.ZF�FkEwo����TU�����e}k�㪻�D"�AX��Q_)�h)���4̘�k���ź�q���S�E����TNdA�MѬ�뫇����O�1 �x~�vV�eI_�c�������op�ͥ������;j
���m�#��R�Ѓ#<����ŲU�[5�����ٝ5d�5^Y��丌���:�i/�2{X�6�*E�8��j�H�Q�O7��	�z?ƶ�O���s:!�'�;���Z���%��5D�{��W�Z-�ͮt)FHX}��~�]_�=�a�xH朆�3�ޙǵ�TJL��f�#���K���6k�6��%%q-Ev�y\���c!�\M�X�7�X3�J�+�9�)�^~y�-�n�w�]0?g��ZU�=��֮���]�Y|��؆(%����q��SRd��T����m���=R��/޻j>� R֝f%��ފU�~�xW*�V����J$�.zpS�����?m����o�_r���F��\U �g�e%�i�&B�8c?w�1�[�����M`z�Z�_�̖U�i�W��P"�K2�0b�42�&�g�V�g3�}wW^�j��D�P���\!ҽnN�M�@�{���O���p(��</K8�nB�.r]���zw��N@�o�H�� �9hi�>��g!Y�]ʻ�����=M����$��@�W�:���7��-UC�&��alm���)�)��+��3?��	zZ�A�׈�����7�LdVҨ"�ۏ`#��'+�h{A{.�2TgX�c�)�8E͝Z]T'_WRR����@qd{K��,��
+-��Z��⸫>�%C-3��Q��:/�\���]kQ�Z�6B9�a�b�A�S$"n�03�^�b3�UU� }%��:g�iˡ�^UE���<�?��zEBߕ����7�#�Bݎ5�wT���m��i��+O|�"��gټ8�T���,�����\���8���r�B�#�c�qW	h����n](g��ج�E7u'~dƨ��f�ԫ#����c�*�����&����vg� Qz�dk�(i�&���F�W�Y�~��x�jo:�訴K�f�������{�m���p���B�k�0o�����{m0��tT�aOH忲�
 ����SK�^�m�1�o�1{:�#�ڔ�Uu��K�˴]68{���CljY�d�m�6�婃�(��.�K��r=����?��R��hAtkx�+�h(_���^�x�|��İ���n ���,|�,V)��'e�`�;$$�)e52��N�S$
5 H���� �U����r@&,��qn���9XT�x�H.� �kX�\NerT��X�xڧ+��t)+����0�ښ���R������h.�c����	P��Ps�}٭'���Z��MlY�v�!2��[ngX2OUKg�sZ��%<�����Y[�䶶z�)�/gkmɦa)[+���(��w݄]�Y��άDe�J��<<����/� y�N�-���V��i��=.��Z�bB�=��&k��a�~���o� ܉>rN��rNDDD��ћ�$�5B�v����D8��dMa��U����Sղ5Y7�vtvB˾����K`�A��:U��FU͖$�4��Ϡ����y	�m��- ��yY�R�<L|<2���~e҈(�a���#�u�1�(�}�j��P�|-I^">"=Wˠ�ZΨJ!I����˻���ɇ	5T�,w|2� .��o��Mֽ垴�T�����}B��c�	(���/tz�0�E�h�|ማ\�ĩ�q���]���4���n�yl.��YtԲ�ԭ����Qq��Q�~���i�t���yMCC�2�v�@�v��Esg�q���_1툻ǘ�8�8:w�4���'2Ͻ=S@��k����,G�Xjrilb�X�JHH����b�!���	�E�Ne�����>g��o���)E,-m��X
�"�9?2	�`��o�<�ϑ��s	(8(O8��yDv����uO>o�"���!�q�T����	�a����X,�Q��\�A�t�K?p�	k��%�s���~:n=��{߈ ;p�F��(��5�U�H�DN��~.-v�Ա���$R�W����d��Q���v��
4��0��b��p�Z*�Չ�z�H�ꅗ��X�`b�7���m�3~: h
� $U�>���)=�H� @M�P�1���wTFANi�U�qӋh��)E��"�,�R����$�R��"'Z�G�kfh|J��.����*ZL���.��C���Ze�1$x"�k��_I:�����X�*�-2:Ldz�Q��y|I QD��T�F������6����];=���"���I��҃&&Dq�S�w��D[��E�����3�a)D�c��!���x��W�_���_P��(|���N5�8��Y�1ч�ŷ�H��M�-�#1ў���fٜ���h��ePq������%	p]�������>a�_"��.E�)>�������v��ˏL]	���*�;�i��l齫,�� ��9���Ppq�����8�}m����I�!�$N
��v��`�y%Ǵ�n)�I��Jr�P`k�B�:�,�gse���))G"˽T���!.�waa��� ��1�U������=���^$!�����G(J�����#�11���a�Ш���,��Ti���{��S�K�uN�{�����-�"s9�yseX�[���*��g!�G5��/^�.��	�KX���g�:+s�p�R�y�f�Ch���G.��qo˩a�*f���v%�x������T�Wsg�~Ѱ��DT�+/�_և�x���K
ێ�N��7l�� �4@g��)��	'U�v����u�k�r���ȟu	3}G�o��<S�X�̑��-T�:�5�</�НA�wmK�����2����J!������+��YkˬU���	5�k�b�~��W�H��h����i��^�a|
B�J�Nk�g�B�[����İ�>���g� Jy�/)u^�����Y�@{���ҙ1����_8��ЄB�b!L��! ����R˃S���Wrni���R'���-�4n�m��|R�xsZ����g~�Ƃf����oC�0��;k��k�4Z�Bi�^sg�p�+1�hcچf��k�Ĝ�3����%?D�xj�u�޲ '�BE���^T�4vt���t������	�,$���7�:���V���N��F��M�_/u���g�Ȳn�d�g��O�b7B�+�4k-�L�%j)ӴR|�]xq����rcs�n=�UF߿��qT�E(3��_Qل_�4��'оƚׅ�ϰ�+�� �<��&��uq�.�8���i����Z�d�J���rn�w�>#��e���7���q{n�OaZw|���6��
5�,O{�F7����KY����OvH��`�X#�~@��#Ŝ�t�f�����oF�emNW��P����� ��M�h�6��|��Y���~ON�֖j|�/����]����=��_@ֳ>B	S��SRX�?�����\97X����E����
��]�9!oVwscb�(�'����R`�ǐǜ��ri���nΊ'D�\/�U�"�0���̲c��v���]��I`��f%4�����/��B�ƾc�d8�rr���V�5/��y<s��t7��h�k�n��ިƗ�9�	 �җ� '/_S$$���`Xu���ܣm�x��ˇIt3���KS���ԩM�s]��❞ans��=s?p��V�q�K��p�45����UW�򯄙R��}�ea�X�\���=~i�Lq�P��ۊ���;�|���p�{��.j~p�]1��Ϳ��A�>��������}п��A�>�������������[�[8�^�j�廻����r|���Hl}\{�6��ֹ��[�����6��It:vJY�4������6�*<����ԎS�<N� ��y"hc�;�'I�0sزn��IHO$�ujx�ߡn�PN�L=��_�*��|[������п?���/yj�a�Ovp2��=�d"|��:�� V�	��\-��4-o�s39�@�lA��c���{��N\Fо�4kI�1Z��h��43'ֿ=�u��a�����.���$G�����Z�2��W�;�W��ǳ���.~��������?���d3D���ݑ��������2���4��gAwm�L��,.P��U���NaQ�=}��|�����Z��}ikk���D���N��E7B���S�����	��o�22����8����69���߳��7����|�d]����qu���F�c�f���h��%Na�Ӄ�gJ2���qv�A������Y�_Fs���2�;..��8>��b��Y���b���J�r�hdtI���=��.�9rz�kS���|�?��Q�t�Ύ�S���іp�"P��x��N�N�(���0�k���>�+>�n}@|���|Qn�;��H���_�������t��[���5>>>Q|�]�?i����w-�$伈�=3��ek�(�X�^��o�S����f�}��������*
�%�II�іpʾ��t瞯a��:m�jjd"7ze�f�2��NH�lOϮ��7�y�j�:7���W��l�� l� z��-5!NA�����Y��ҹ��ϔ�#�5�I��Ų0dHa�=�D7�۝��~��}{}�����HG t���Id����W%/�������W��ȉ��x@�.�H�9��*A���>�bܡ�Р�h1#�Ց�/[���u�Z�}���"M^��n]�Þb���2���&�,������D�V�.AS= ��Ȅ������PC�#n{���Q��X��7ccc|�{��5l��y��>))I���LI`����}��cIΒ����"R��
�-%�P�����ֳ��Qh��khh��v���_7SRPxc�������d]]�a|�s����i�/Ow����Y|�?�U�/C�䴺�v�Ft�U����R�<M?���K��>�7��>��o���N'�b����`+ 4��͉�^��G �� ��\ǻ>q�Uy��Ub�x`;O��R]6�&���u����b[W�Iϥ���ozA�����;�Q���6$=����~[��[UM�---��3�@!��ѩ�a8�_����#B��҃|g�:��K�?��Q��w�v�n791k��ds���_����0�W�����,�;���g�_8̢v���.�9��uNn�u����V�%���n����kx�}���4
B����f�P[�nw�����E2B��E��0��������K@����|�zG�[o�X����t^۩.�g~�����f�J�Y���	?��L����y+P���@��K���e�3�~q�O�a~�6������nP#[�)����G-�`���=S��n��7�*����yY/NǾ}�ّlΫ͑�11�)�WD�]B�toJ��=�������������p�L���>�i�`?��-nu��n`+�(!�O�i�Ĝ�kH4�TTTgH�̻��M}�N���a�.�de���'���Ϫ���޲Ϡ(���4��/?[��ڳ���<�e�F�;�[�}��9A���+.H�8"���Eo��҅��Q*��K����	�q��a�Ӑ3��4U��&{JD��4h��(���D��[��耇�#���ď����g�,in(
��X'Ȇ�8�L���߭-���7��#��io-l��9�-{�ЃZ(� �nc�'�� ��Av,�wUT��S2�l�eA
jj�����A�(<�d�b�b�u�����H�uP���GI*�����Փ�2[8���4�������	 L�(Jݐ�����Քr�_㩀u��q�B��>����򚵘��!��8܋OAW�#�h����#�ݾ�f�yg�K��\]]E/���gb>}����5���1�����ef�H�½��[�6�a��% 0�Sϳx�\��l%e���i��k֣���n���h�[wG�Z���CRZU��Aqѣ�A�;.�-���������u�����
�%�fm�������=���>��:w�����-��Wr�����-༅�`t6�W�jd�L���T�ڵ<S���F�Bl�,��r������luq<�Wr%�g��M����3�?����$�<L�=V��I�;���a�*�c����ٹjέ��J_����ȜK������P�y;���(, 2���맒����)�P��X}0�y��R�����MkJԛ�N3Ϙj�Z���د!��B���ľ�<��t�(#G܂��dϦ�G�Ŝ�Ue�]2�����玴�9�����x���U���RT���D:L���z E�&�5|�#p{eEE��I(��b\༱JX�p��2��(��N�ohjj�x?òC���&G �魍[�@됈�4߄1T  ���{!�ްR�N雤������i-��w>f)+�� ��L� ��ut��V^ԭ�"J]���g�?�[f�a>/&)����DJBٍ���i��r�����VpɆ�r��w�����`&��V��pAOo��+�V�Ü�C-��۪������E��i)߾=t%m�cKC�:it,�"�>Q?��";,Y9�u9d�]`�	����`J��Ւ��a2��O�\	ii���9���Y�I�	�)����e77��}׼��#a�k�Q��E�c�r\'�2���E�v�{�����xI֪X3�`J܃��ۼG)%���]�%_kCCC-CA"���Sޠұ���UNS����p/���r�n4	�FS:1�x�fmdd�uq���?�Y���l�ΎZO�����D��z;ভ��s>��ʳ\k:�����O��´��ևN��"���x��4z�
ps:\��@1�y7{)7O컄�|@��:=�s�}t���&�5����*:::��d:�贠@����
=
��,�xC�G?�`|�הx�T�����OV6y��m�0�����v�-
���A:3[=[w���S�pO��� �b����M����RA�	�e���|q�_L'#�J���GyM5g�	<7"�f�(+'?�0J�пR���SȊ��PZt���S�AZ��DP����o��@�{����jV||�S|y��ڪh��쓝a��I��3ǁQCh���������W��������[��L�Q�#\jmk�=�@����t���O�s��W�ߟ,E���9�P��O���w��W+CE��ʝP%�	�=�ಚ��"BC]�?�`��2�C�'l״sĮ��o��J|�ي8줸�.3�4,�w��88|�ANJa��iTfv�est����"�*�όv3���S��b'yg�ǁ+�ĸ��r�۳&�x|���ԁB�v������'SX~ܷͭ_W���b��=ǣ�J�+}G�g(������qd���k��3��k�`�0>8iu!����D;e��&��x���C�(�����}�=+��{���QyJ�#�n+
'5���èP�6G�Ό]8fm���a���C}�+'ZoKċOʘ6�?z1**x�)
��n��2�/��EN���a������� �D�]`e���v�EK�8�E��s�[�e=Vͷ�F�7��$& z����,�EE��:�Z��-%%%�����견�ϫ��_/��,a?I.ݚ���h�<T�7������Tx�5OZ*�F��ucF���'''KVD~R�F5��	�y����G��M�C)��oNK��������*V�Jt�����}�_)�g��x��!\Z�i����9����1��Cp�>�{�]��6AO���ɯ3�#L f��P�թР����=j6���r�g���{_O����:MTRB�����M�K4�|
QB����(R�2�2��<��"S��Sl�m��w�]t��||?����Ogx�}?��ֵ�5�kEiv��YY[[��������"�,���!����S�8RZ�/"u��"'[&��&����x�6N�.0m�ඡXid�U!�Z��� ��ԅ�<����p��3��V���Rg�֛D��03D����hG���N�rҖP9����]i����!!�N�y��e%E�6U�O؉]X��hŃ�-��iZX�<X.�]��;rywz�Ǘ�ja)���آ�>���H2���'��
�t]A��oߞVk-\�� v������S�BKk�yt��Ӽ��R�*}C������{͆c.��L��-+3mO�~�-i����U�CD���ȧax*W�ć�(mp�˯m�6+a&1�m#����\Q�C�ⲱ�@�Z�v^@���M����x��n�y@!�,y�6�_[O��n�S��9�����AK��֎"NM�w�����S�˺:Ѹ��<r�G��9׬I4�쬼���j;v���a8�B���!��q�����Z�f9��2?����.�߄O	S^�v���p.\`���v��e��㋰2?��j/1�C0蜆���5�}F|�f�	8�WO�&w�/���Q��*��?�CCC�Vsss�t���xU'���W������Ը��?a� �#��o:���qgr�	vZ�|V�����4�����gS �Z��?I�bF?۩��;>��W@�Q���9.�n���1���)�G���N<��b��[��,���p�[�2����v�̟��ۖ9���"��˷xd����(�V!�M�سg��CS8Ypt>��F�ovɢ�RH�M�e	�	k_��Q�PWڱ6;�v#�o�C�-���Dܴo��>�Ɵ�t��jI���΃�6|�|g�Y1�!e5ܫ�Ď
�a��Hb��ƧX��%��%\�i�J�F������%�+_�l	��
\1���u����CC���Z�5�2�Ǳ�f.�Kd��a�R��m*_�]�Cɜ�E1�
��uI��G�7/����PLl���Lǈ&8��
��>�

�}����Z�r��]�ZȟJn�<&--�� ,�l=:(-�s�cnn����8����p`��l�>�xDw/O5�����bɞ�=�'l?��Pw~���P �yۥ�f����"a�
M��INz�Y�r�r�N9
/
��7����׬�>H���;���N���Q��z_ޜg�}r�-??���03,�~���jex��9��kE��-�\�y��3���n�L��+�$՟|FG�G��/}�>3�;ut&�3�������W�����T� V��7�[.˷����~�&�_�(,�#^� �t��2	�u��S�ԟ�ߤcQ�;D�ҷ
����u_E�)K�	*�N�����xg���u���ԥ��܌�䕦�'�;cʰ����\w�d�I|ǀ%H�Ɓ�2sj)�ئ>0p���xc]�٭�5{n\�+�׉Z��;?�?5U�:�t���lŗ�~���z�=�5�2L/qK�C�����2��� �aaB'�I�=8�����_hF��u�5[�e����s)�x��>W� �_��8�K�?*j��M��.�(
54����~/66�N���u59D5���\Q�/��\��eZ�7��CBNY�� V���ՙ�88?߬5г�lA/�_�����H8Z������S����N���l�M�����HZ�e�:��^_[�e0�Y����/�%�T��g~�mo�c���&����ݞ�3�x��}�1z'm����CҤ���	�}��G�i�7h"�l{�ͮA��>77`8s����/��= �N�|�+�Vk��^5�S��Y���JJL�=H��T��%��RK�2O�Ht��v,e����~�xƧ(�����խ�^�%�G��}��uǷp��)��C���?��7b0x�c�ZQYy��U�q#^�	��O<״ܾ6N_���Lb�|��x��d�J3ϣi���\��,��0�{x�T���V�s���Ǉr�5����G�cfYi�Quuu�(�Vr)���������aa.@�ŵ*cue�T��G|��ˏ;5������߿��SMz��MFS- ��5�D�=��br*p�B��e�ڷ��R�6O�@�L���MN������}]���=�7�O�bb�2���y��d[�c�����Џ;;.X��Bу~I��r-�k�dݮF��!k~!ޑ�h�@�{tJ���t�G���LQ�/��<Ϻ�H7�]1��踸 �
To���zz.8V6���[s�H���#��T�هSi��\L+>ԣ;����#aaWp��LQR`��k��ʂ�����G��'�tdV|nD��!��q�#�[N?}�����ѽJ^�m����?˱��X7�߼�I�o�b���	�b^p�O?���NPn5��K����u�e��}���4�<g�j�)��u=>t�,)qww�r���_6mO�QY0���Z��ΐ-�c���*1[�a!��]�Q迫W snڗ�$ˉ��S��ՙ�$i���}������b8j=s��0��I���+�1���f.��<�]-�Q��r��Q1/��z��u�8dii�we��>�0E�G�p��&h`O�iJH�慗r�y�{�n��d% w��%�2�q��Λ�tuu�Z��'߂�.���������5:!�9���L���3�5�����y�@J��o�W��m�Օ��J}��e���X%q�k�E̟d�-��J*��j���"U�խ�[�	�Oc6�����6;-���÷1H���h��UO�i�ޒkk��	V`���B��n�L٘���1��^^��z_&�bB^II)c����D�9N�|��j��ʡ��#Kf����u�ۈa�R@�F�<�r�8RQ6#��=���cKsѓ,����m:5��4��d����w��S@&��5eOV;g��3�*����j��/y�j��:�!
�H��Ha�3g��8"nl)^<	�α����u�<�J����>��-@TzƻI�e�4%3/�-�-k91�#�),�7`��">jƛ�Ŝ{DE);�d=<��Q�	{��P�K�R�����ۓ�k8����z�U^(9�����~��_p�VK��=1[�ݷo_��8=U���0fS6�汹f����cbz�3͊�~]5s���S�R��U8'��9T%I��3�e���F�oYU���q�P�y�"�,vj��Fx}�#M��ߊv}aٓ����|���N�`W5lƆ��b��.e?��]�)�%C)�YuO_Gg�J_C��9��K���(LxaCaP�?f�������;=�G�HB��{�v'��b7Y�۞��Ⱳ���w (�T�mk��pӾ�H�a�H��#�SI�s���[��0�3d��f�#{���YE&0�xoP�KRW����mr��7F�����5���|��G�h=�3�OtE��e����)�d+��&N����wXG�70����M�c���UU�y��曰�&�9�KQ��mXp�BU��p����;�+��W�G�En73��@W'��f-��>2��֖�~$+�j�#�d4Hp�lI-U��
�x�-�☵�Ϧ��g�a8���fM�J�v���L{�k�UW�	vvv��PŘ�Z����H�D���8�+0���I��z��bk"�o�'�%)=���ji٢�Y��,:&f�8*q��<0d�x���8q������;3z`r���:�����ç����{�S��>�N,��&��a��e3F"��K9�8/�Ő�C@aE�LkN��m���� ��	g�������\�-\vD�uxx�`B�ߤ�ƞJ��O�H?1�3�ăX��*�6���M&ld�tq��K8��_����0�H�P/�߆�78�~���oW��s�F����΂/�}p����ؓ��2NxԢ���^p���X���D{T�p�7��X6�l4�6��-���o�
y��>j�n.64�k3f�D��\�V{1Ք�����ʀH�U'���*3!Me�mw�ܪK��K���|�ʚ��S�=�Ŝ'�}l��R�UR:���cR���2�H��ڣXIbr��Gx�W��<�\��䀥s�3�S�Ҙ�a�G4�=q�%脏}�S(F쪇UQ�3�W{��1φ�;S���6S��N�i��^�4�N��g)��(�����G�`��t��KYW<��QUDz,1�WnIJj�$M���E������ݠ��5O&L�p"����
����bҹE�u���'N��$�\�[�b2I'�-�LQ
�^ge���p��s��V\�av�!*	Q�4�Eb��2O5Ota^#c�`W5'��R,���6z���rK6�G�߱h涍HN��.��� �g@��f�����Q�d�����f@>�M��2E�Q�z"����#6���Z�03�B�t� �~�����Ѧ�B�	.�R<��DNa�򓗨��9Z�r5K�k�L)��p��њ��@O����8V�	�Z���S�GYa/5��1v��ɺ-��} ����෮�ȫ,�C#t��ZtQSDOܦ�^	��c���{��N�rqJ:ޟ��ȴg2hoiq�;����/��dn��Ln�bt�,y�%�s�e�NN'gV���M�q`�v�YUU��,ͨS<���Br-�	8aCCm�Ί���8l��: `	��|*N��e����ʌ^̫wnTz|CG'�l���$j`��q��I/M��b����!�{�W`�a� �U'�+�r^�g+�R�9.?Eq��LشTAKӭ�Tqt<N�]��u8�$��N����;މ�'������@l5����&�{Av���.�z�-<�s	�`�����c/9�G�=�V�R��.u�p��F}��h�X�k�lVo����p�N)���q�����:_V�o(��|h�\��ZN��p\�:�y��2��i��9ܦU,M�m����f܃����i�a�<{�*�]�}���A��B�'Ombg��ˠ/ee�&����Ȫկ�����T�h�cReZk�}.�K<�H�=�%����-T���+0��8��q�؛
z�4�;���c.\�g�ȈД��h�	�!=���	���"�{���3���Y�y'�Ө�L������)����ުm��7�їx�>�i�T)�y�š��/9p�)}h ��i:��U�w��;Q��}�V��Q��(��AHAA���'���ݣ\,����PD���1�J(Ϟ���*�D�鴯��d�K欿�t�	��^>m��%���������fg�I����roBC�T���ʟ;��H���Zb���2�5�6CIXh���l�s����H��'���f�E����`X����Zp,��΂�"����_Q�/-xx���<C�l�������#���Tb����e8��/�g=�����Y�N�
�s'[m,k'sj|�_,�?9i������?V,^\����^g�F:�?໽x��3���v�ri�\pA�t��خ���7��x����˥j3$=.8�"�Ʈ�T����;�;���_4~�x�\�ְ+a�X�x�h�3j��k`�l
q ���x������ϊ�U��E]V����yBIo�í�41�916�}���5y�q��?�K(�dei�Q�]y$0p7�ͧ��_VF��7+?$8XQ#=r����њX]��]_�����E����g|VRT�<??�a8�%\{�O�$@l��;�YQ�8��=�Y*h��好W1�^c_��������.aWt�^|�e���oਧ�o����o��w+�Џ�k)����@��g��"C]�3�ht*3���������ɦԧ%5���g�(`���
_�:��a�&׷�i8������wY��Z��Ml�v�H�S����2,<>��o�煽µ��m�\6�k�~H�|�$y.)q�;��HKKw��6Mx��A�
ݒg�"�(|V#�M.�	�M��u��z�Sء}�	%S$��%,E�Ǣ��0����
Î�ab����_/b�e�@`G555�ļD�]R,�4a�������N7����e�A����W$R5T��Y�]i8��Qخ?�m�va 6.q혎�H�?6��i�Wv%��a�h��{<�N�*��ݭK�+������eVI���@>1�;���Mp_�<�#�����jz=�X�D��_Z���f�
�p��G�u��pj���}p)�6?��Z�����l��.��������X�|�c��E����.k$���Ǝ�فW�6��b�}d���u0K�݊�H�2�*O�t=q���A�6�mń!H�ʇd��:"rf&:l{�em�G�'l���W"��v7��B��l�%M���CX��g�2����֏W�U'���Q|4a-ࠠJ���=���Q1���v��2z�����{V� C��"��I��]ٱ4��-`h�^��%H���	��P�8�W��U�zm~�E��Gkʷo�8ph⺾��LHjBkg��sK�y�K��R�o�\L�k�]C�[�|�=C�U�l8�ߺk��%>y���}�Z_����iǬ �y��#�s��1�:�1C�Q�U�0rZE��þp2�4�#`2�>�D�ޒ�NZћ���v@�둙�)oWC�Y���>��5�������5:��ص�^��Q��L��k�ʖٮ���U�s�e��\�24��\�`�w�|n���닳k0�=���#�����%�R
|��C�~L�������ȃ�"�1Ow�E�f_(i9x�$`�ڊ;��=@Y#�8Ï-��1��ʗ@�.�k����R�Jl�e���,�6<����
��39�ё�J�š�G-ʐ>R�2X�mԢ�m܀4^�o)N� "9Y��?^�fٝ"J��u��i~+��qXŹ�{�?�8_����a߿��&9vk���㴗H�C1��c�s����~C��������ӎ�������� E�jVg)���^��r��X�I�k� �]��� X�U8��E@!r���:�^���$p��ޱ?ו5���
֌��e�c����x�Ӽ��<4_��t<�,mμC_�c�a1O���>5������{S��w�C��?�m��U`�C��A�S����y���c��n4Ύ�~ɇ97t�%#\�=�T�@�81��G)\8,��}�T%v)`Hˉ�?�P�ׯ_/�y�/9��t���_rG��ֹ���dԉC^�ԇ{�2����d	v�/)������͛�����pwƵq�0��������=8P��е���X���!�ԋU����,$�ֈܼ��=�X�7U���M��9'!�,tm�q���l:8�*������S�Gc[�F� +F��m�h�|���5-�'h� �F�rCl;��՜�K��	���VQ�ʆ;��}�S��|V���qVI�J#��[u��Y6=�d'v�޲�m_���u��Җ������R��1'��."*�%K5�k�,��H9j�O���	����>����m���V�kp"5��kĩ�X�����.�O�V��x�������:�W��8��),	��>�ӣ�`Mt7PeɚЌ��= �k����Z����Сc�<�c�q�Y�*q�/]����=Y%�q�9��a�IY����2�ܪ�hüK>�̯ͪ��Ф����K�2����)����ZD�_��5v �X"�8ʼY'x�ܸ����Q���)��x���P.nf�i-�F�R�Lv7�Q��[�H���w���Se ��Z�I1.f�]f^��t�ȕW��[����x�w��e$_�r�Zm��T��y��8c/\E9��&���]��Mȗ�ook���P���c,hG�}�ὔ.=�Ӎ�S�{o7�uE��8�sBcָ�I�bt�5�	���6�0#����$�1o3>PF�ݣ����o�놖On�.q,����5oa������n��(�����Bw��L���]6l=~3�E�U1��a���삊�h��Đ7�����k�pK�V��7�`���Y���pn"�p���^1������Z%��ի�|guuC�Gj�!��'J`����4�:N����a�|�ZG���$0+�8�u팷IǋZ^r|�I�� ��D�8�
�
/�ڎ�2����=L�$�_����p�
Ҋ�x��c�^���� ��{w0���{�&{(��-�����Q4:��
4hmZ��#,��J���2N��w����§횵�ۿ���?{�H�qŰ�Ga����0(�+G�"FFF�JX�����+��+�)j�1`���GV�]=ι�!3��0�h�Y�|<
wE`�璟?_3;�(rv*�l�p�}+������f�!>Ak�
��X�%�.\�������]*�gHƙ�xR'��>q���V��9��ۆc��60�yc�e�In{�h�N�RG���	��{Q$2]���9��b��"����ɉ!��u0OPI&�L>:������J(�ꧧ;��K���_TF�s��P�^���Y��,��m�����#���bpH�؄67<<����	� ���r�Njc�g.T�kJ˵�P���[v(<��vDl*$M��[��
f����Q���Ka�É��"#w�=o�`��_gU�]�
�:O�Q�x�Á�,�k�ge#&��UD_��d~.�]���z�Z�+*��$OO�$�}���S;IY��nO�a���I�<R�6xM�΃�I뢫��p�И�vWuԠTs��צ��9:ޫ\�ϡ���T��E�gX(F��PMޛ�Æ��qy7�y`Y�Z�M��,�霮S���VHZ��#�u��V�a���={��v=ݾg�k��?&�m�u%a��2AK٢5e��h�V��1�|V5��oc��i߳�,6�h�3y�DX1:K��˟��G����hU��KE��b����]V�U�zU��Ah~�p6�If�)�ŊGY�:d�Y�x�Z��6mb|�}g�Y�Qm��H;ӳ']�M�"""�[|�,��/���|�(�7T3�����a<��5��#���$Y��^�&���wj��[Q���4�y44�˹pע^Np��"��!9��]b�5qM�|����D-Ak)���h��Dtg[G�)��pv�ޟ�6Ѥv��ɫ��րR�糘b��,F���JIN�����4:4�}#@o����p��^8xw'���x� ��Jϰt$
�X���U,?{(�:�?�-�cl�g�ཌu}7nܘmY+��Z�B�5�)����Qg���/a�� 
��N�O<�,����ǅK������<�>CF��MO���q��C���<V�\:"� ��c�pޛ�ڣ>*�驸�ӫ6 �׾w5�����ˬ6x{��0�f���=��"Pa����.�c&P=5lZ�7��j߶���e� �Rk��;5O~�$�`�zF26��\e/#;��ٺ��j-8�M�� 8ʶC,��=5ξ�k����˸�.G�d�Du���+`��A!8f�x�����,3W�=e�����0�/�<�>��0�xщ�j�6Z�p-`�>�D�N]��S:�Z�D��c߹E�>�#s���n�Lذ�J}��G⣯������umm�2|��߹bj��c��q���E����
�*�r�~)kd��N�&�R�D�ׯ��V�$}������7>u��E�Dc��H0�,[d|�J�X��s�������_
��Վ��^0�8��l��ݥ:}�4��U+�k�L��]�6�li5:���/vX�
;�`wkV,[w:Ϩ�x�p�.|�S���<���������q7��3�������b[2Lo�!v�����w�vV�����b�R�+�>��� �3U��v�j�p���"]<e9�p8�~J�� �Zᬟ.p�?IZ"��:��S���z�GDWq]^��E& �@�]9E��ZW�ŚH��ĺY���i�n�C�ʧ}�X'���3�p�N�4�6���=�*bt���2��b_�Y���^ت�����<�>~�����)�>W��@�j��|/�h]�6��.�6���L��@���ص&�s+�]��9>�7����hҢ2UK]�K�#�����F�!�.��"fې!n[�D�0i��,�%������w=�I���>��|���@_�1B
��,5�<}�x�Z�M�q�רW��=tV�
�ձ iΙ2�vn�g�EC�l�Vd��΂��~m�U�.�ʲ`Pjs̍��`��K�:�Y���án�;�v�Z�o��>S.�E�.N38᫦���ʇ�:�OjBZ�:��΂|E�)��-����m,�ĆjI$3�1�$z#PQCia
�GS��� ��B&f	~sT�)��hi�G.�L~�����4p�5�a���%˿~��MK�OՌw�Xez6��A/�-и�8�%??�\b�CI�_C�7�T�ǁr��E��,�ߤ���i�A���Ö+,O �����������d�4�,X�Q��:��bx�M�
}U>�e-'�6�G�!ٮ���a�N
,�;+���g��s���L���za��FR�nT�u��e7q����Ӏ��ᓹD�ͯ߸��OG+����,�,�VO
��tJ�
���CH�LjڻXzi�%��� �Q�#L��i:
��s��X��w�i�c ��#��D�������'�?���
�$�֣l;�cc/�*�}�t�I{!��G|�H�c��ަ<3rp@����Ւ��J��S7�g�}{���oz�C)�Θ����Wֹq,��Z�)#���QU�1���-b�b�ir#��[u釮qｵ6镓	NG�cBZ��)[����G�nW�ƭ�)�k�K�z���fP���@1~n�
+��G�9�)�@C�#�W�:��V��`bp(����Y��`nƝ���F@��!��088�ea*�X���G���켢?�0.�&�]�E�8�z��_q`Dop�J��t�eb9v���V�)^�w�ܟ�%2>�M4��|Y�w�����N�]�� ag�u}������@���5�F%gz
LS���I��3G=���l  �9D>�Fˑ���F���wE����+w���e/�>� �$�H���S6�Mp�i�=
*�b|1l5�؃�6����ΒV �R�ۻ�陖/� #�0^�WFD�U+�I�	�W	0��gs�t:����A�HH�#�����;�`���g�#�0��6(p~È�?���R�jc�����q���[ E��<�s&r�"YO����������4gT$?�&�� �m����ġ��F��M�4P'�P�'9���ݢ���v�+����|����Z�}�h5C��8 �i��qz6��`?S�w���>�1�/_��ک�I$�F�P��̚
��������O�_�~��h���!U�x�5�Z��6aN,�2/۱A��	J3V%u%���t,�4e�|���&k_�?;����Z�w��%i��'���̲��w ��"
|�Fx7���@���4؊��@>rʢī�=��3�jKUtk�ij��\��`�����5����{�:���J��]\��5-��q>��+c��yu�+w'c��,G� �����t`3�ВL{������c���k��4�5��-7�!����qd�;�C�ϟǌ��V�[68�$Hj����R�����3�!�+�{��>^�I��+e���O�LLܷ���d����L(6�*��ldz���{�~��YY����x
o޾}��n`�q�̒2��`ߐ��n}�� !)<�ϡ:�����qO���{1�$�`��] ��OJM����M*xu�u!4�F���+a���[�O)�]f_�T�_��q�?�����(�|�[�4I��St/��Mw@ g3��+q�M�yByv��,O��!K�ط\���[cÇM��]�q��V!�	�eimO��@?i��0��$X�V �R�d<�=���%�P��2�]���Ko�:��DG�?[����]�8�#Iv\���C��
��'[;ʣz|���T�`]��Å���ߜĮA7�ۃ�[�Sf�)�{���.Y�sc�3V�q�3z�����.�ݠ��<H�7[z*:�����:f��wAE:�����ů��B*����^�J�HMUU�����F,g�jXIv ��(o;�UV�xp��[Ш�{�7	�<K	 Vl1ر��<�>�89y���fM�9�M��o4>`����������(/�v��浙Gw��4�]������իW��C7����0T�H��a�jvl���I0�$�_�6���ý�cM�Zn��"��w�N9�>��_Av)�an�:r[q*��C�B/G�Ǹ�X�z�}j�o��K�4A0��_8%]�̽��i�	�NN+�'�:Vq�����R�Ϯ9�`H����sI��.q*��k��*���tC[{�MmWu�uo�2n�B�zfV�_[br�a��t�`��$�N;z�9}G���H�-�P�`��$�jH�a��a��s$ǒ4�w����
ޓ��%�T��q
LD\�4�t�
� ����3��6��a�Pw�KYYv�x~��}�w����3+B�&N�Ôd�`��E{�jժb_�Ѳ��I����4���߷��ֱ+8-�4�]�>?�7��9����7M�����.+J��8��O ���#m!+�?���ҵ�;9��Z��cv�q��1�|���G���r䐞�c�1�ъ���7����S���{��?HUhUq^�+є7�1�����|��;8m劁��2�F]N2�}��?vc�|��wv�"����T�[��W�GT4Ǖ4ֈ@��i�d1�b�r�����h���8���)U��=ZC9��h������=Y����d+.���*Kc-Q�:ǃ�p�Q���� �|��6�����*��j읉�1��LNO�,�
����JO����ug�+�p@�x�={���
9L��?�2s�ѷ8K��VI4�7��Q�`.��c$�8�=�=H��D�}�I��u���z�e��t��JR�d�;X�c�aGo�?��w���	}�pV6�p���"zY���!�]��.��y�ڱH�<���آ��K�.���>�'5i�L@���h%����̙3�l�/�)�C	�
�>���̂� ���d��@cp	�ᳲ ��˴@���m�� 4�	C�3mqz֖_�������=X/�}O��e��'2��5�'�/ *��-Wp��L��a��s�?�ga"�O)N��-`;��oo���8s�KX�'���M�%oaJd_g�;��j��u5wg�U���x�}�YJ2�>�[��]�IWU�YW�;m�'�]�x���I�����uAӍ-&����X�7����c��?�:ꊭ�c��	k�M̖��]&�R���+�477g���}3S�k7M5ei�������
��w�FJ���O��1�?1Ү����������#5p�lk��n��9dy�S��KN�����W���7���Ͳ��[���c:=-�����`�ã:�Cd) �a��;2�SI[;�����Z�w����B�e�#���L�͂��r8�'w[�����-8Ig�1iC�ëAij	/(8��R�1�w������*yZ��b��;t~�76N�܇E�F���9	\�#8�68�-�ㇴ�a���om��]v����n$���Jp�����cSE/V���(J���d{U@��t3�^�%��W�K���fF��*<�
����Z���dsێ�F��c�6��T�F�S_-�s��gރH��K��w��z[������L��v�e~���s~h�N�J�t�MD��"�3���m�����G��Q�dN7�����d�Ν���qbV�n�sT������mv;��ϟg����?�����3���?�����3���?�����3���?�����3�����?s�R�\Vpg)i��D�����2o����rm�x	U��|Y�>�ﲻ�Ui<^��_�7�7qw������Ҫ����{���̥sΙ������kϙ�9�;<�ȂD�d�%���-�Bw�]�t-JTB�H��<GY������b���w��n��K>m*�y�]s���1�����֒ �$��S�>u*��C�e�F*C�5�*uߖ��&���v�Hp�cIk?i�����G���]C�y���V��<n������>��o=�ݜg�0��1�=q/ײ���T��ظ�c�2�C�@�[�L���o��R)�PmP�}a�c��MrQ���2����~�I���n��D�ge�����&��,�c�K�=�"��]��F��fm�/���q�,)`#�����&�Nq�yyy���ݻ,��O����Ax\c����{h&)l����QS!�����ptib��!��b3�\3S�ď^�Xl\�E�NQտB

�����Hέͩ�s5���pk�{+��.��I?�,$롹��J�?�*�4vޯ��Fv>�{�z�#M.,,�q�~>�}�3�]�����^�)R�> Z��h�m����2����Q8&?�u�=\Se���p<�$�g�Y4m���#&:u�f�����7[���zz{W�&
��􆧍w�ON`IV�� ��1gxj����2H�#�NN��"뤶D��D�q�7�%�����{V���&ܰ���HT��İQ�W�'Zu��%t6�����`U��N��x�D�&ovE�?��W	
�X��*-{ėB��YG���_]��9qK��	��~&�=�܅q���_�8�2g��v�%W����~bN(T����A�Az�<�dY�(�!��D��Z�dp?R�����
�;ȅ�1�)#7	�֫ch�u���0'����9�����J��)��V~Ӌ�-γ��zQ*s���%�b�[��q�H�y�i
�9�>�Q�]#���X%@�������M��c~�k.^�
��ʲHq���zM�PFI�y��vV�:	���oFxN�_��G�%�;s�,������f���%�עn�x��ޫ�C��j�$s�bJ='z�VT�^㭽Gڎ�˲J���W����Q������/o'�� =Ir΍G��Y�]O_h"Σ�T}�2�-2���^��_�\�}�w�C�MKʪ�"Mp��:�9n��/�ǁH���$La��B
���y�f����ؓo�&(7�s�e���tC1�H_X�{����-Q�څ��ۭ	�ⓤ,�36�U־G.NYH=��M7F�75���b̭R&��+���w�.N;w�j��ŋ���G�`A8�,p�ݚ�׷k�,�������R襈��5	w����Ȣl�Y"�[���QP�/�ע��q�TH^H���KZ��2MU���BM���4��n���g?>G�e�j��ǭ7��i��W�)J��_�8t�h�+#��Z�Kq���V���G)tK�1㢃uO�����kq=@��*`9��~`=|)�7��|���z"(b��b�U�*H-ǒ"\�]h���0<,V�����}5�4t��.*�����rs �ƞ��;	k9�wl���٠��F��󯭼��Vr���Ee/~\BN�zc�S�z3�$��_T�������	M�B���"N������pn�!�����nx��cue��c�%2j�@��kz�I�/s�����)q��?n��L����>�3�V��𮰘�ӄj�N'����G�i��O�S���$I �x������¾�<B��H��ǸoX�R�E6+n�3�����q�t��[�x�:����Sg�m��$���&��Qߴ�Z/Oe~��IxHO��<�ll\ 5�(	y"�E֍�m�~:a��y}�~�|����2�@d�o�������h'�E�/��B��k�â]��׾k��Ѝ�^�쒒�&Iq�u0�Z�F>���-B5\};�C�\S��h_��?R i�5�n�p'��ՙ�<}�ݎ`,��o%m����o��7�㿝���8�\@��@2� �8�6��wVNhc�j�5�����@C�����������6K�g��������_�8���t��e��.i�M�!�u�� c 0ջb�CH�x+��Pǫ��%6�@�`�G�|鴣P��ANc]��R�u9�8�I�>�;*���	�edΐ��
 �'���E)5��c�$9Q�e����������_s����:��W����,pX:^� �'J�ZA��I>�R�����~��e�z����N��-��ö�Aן��Z@1���kQ���v�b��婺������0`a��X�H�j��گ��\���Q3G��;�D_�09�i���ђݿ�)���D����?=.�:t�����DF���i)PvQC9zd������Ϳ�b�(Q���RŅ�^D"{�N���-t���(xM)����څoE���5]�3<��"�4�pH��I�Pa�6XE+"9��m2u�tj��8���%��/VgRQ
xtu�D���
Xc��N<{�
w���p��iX7�up��J��+�@�'6?Hk(�i}G&��w���j�e���^�UR�1=�'!^��ΜA��>�0�WG��ve�E�]s@���D�H�%��t�i�>�9C<�>�:OB��\@�\T��R�!�
�ө��_�&
t�W����wW��d�u���`�,���ٞ� �6 �3�BT�Z�������5��v�9I��g�/�:%���U]���q[���g��Q���D��F����	'���|��bu7hZ���1$kO�V�&I�tHv>
���^du�k�o�����k��,'J�H�B����b<�`��q.Y �~z�c۸�S���E�vW�u�]�gzQ��z�n���k���]s5^�q�c�*��n|Z����-�W�����Q�x4FW!��ȭ�%E����
S���pO�Zu� MrA���e��� I�ʄ��ӸiI����)�a'����;@��{�t~�����ė�-&҂1�X]:-tK���BZV9�J�#�vќ� :�{4<���C�L�x���2�շ�>������V4L� ��8;�)�Q�}*3>��9c� Mr	9R �j���V���"D����\)46����[�DK�y��_p0=B�jd�8SK���6�<�f�"��}�<�+�p5��z�8�mٍ=�Iq��}���淏2�W[�7�� ��g`��UD�޴�/0�Ь���#�(�"֭j�W�T͎
�Zi���D���ձ9ei�%�� 6���Y��ܼy�1��*c�1�=^�����3��D{��^�axh* ���'��!��e��z�==;�_�q���	'r���;b�p�㏛�)��:D����T���YWY���Cd��%w�]��/櫋!|�@�n�&.�z8��H�8��K]n�I���Kű��v�v�$����f��vuje���(���AZ�9��5	�g��a!���M'p-��%�����J�G�Ѫ+m&��[���%�k�wl�btu���)�qYy�L$&��~#���������O�5�3s�W-�M���޻M?�v\���HD
/��>0�.�ۙ�x���Mt:��ӳ�h����ڕN&�B�_Q!���y��D��	[~*����Aʗh%���^N��,h����+����#n�m���_(I�4{�b�U�AXhû�{�XS��a��B[2!�1}�4�m���Iļ�+���0���@ǒs�Ĉd��
˸x�6�a�?�"ݓP\V�0�𮢢�s�����t��1��0��"�;v|�)X�[C�-����R7���<�+P����:ό�p1� �ʌ�����J ޶� �X�:Zp�8��	���Am^i�1���8ö;��Ln�%�p�]rԑ{t�T`>F$�U��rv�	��F1���1��&�t�	0to�[�V��U#[�N0��4=
.n� ��y��X�؏0�?�ឣL�C�僣dV[����c����'��t�
��-��&�{p��,��H?uNN�LiT&���T�\
��a�t\�׮�՚��8Q��s6����a�4�G H��:Q���.������}����Q����G0�k�p�ȕV}2e�1�
T��3�&�|-����<8���H�7��FÉ6�a��i�TѼp'���~���n��8��F,���ӛ��?2�$7���G�G�+A�(�;�D�r@�$I�r��	��7ږ�!Ј�x�"YY=ൡ������6Dr�u?���J�UND(mȋd�Y@$V�@Xf������)�|ȗX]X�)VI̠�!��~���~��ϏW��N��PE�TB^�7R�^I$,����_�Q�B�pf�cX{�83Q̥.�{ٽ��#+���D�I���w�H�&Z���o�p�(�d�W�t������A���f/�:��%��xyy��m��vQ�V�v5�Q{�W h�D9���_NS�9O\\�����r��9�yX{���J� �� ��XWHdӭ0B ��F3����ɩr�0����N!\��X]�E��捱�;+��c�� ���B
�����2��7����-FƟ�5��{�&�����Q��k����W�])�����U��D�����S"��\K)�,��&ft���OJJ�[@S�ݶtꛏ�Ѓ��=��mi�	|z�5�7:>������,ߴ`2_���tC";: 9w�F��7:nz���᷏3�.��y\`���2��Q��P�ħ�`K@U;��-�����MO�����2���M6O��I�0Q�,�ۿ���!�/��$��K�}�����]<��/��0ڗ���a,0Q`��5~3�@R����4֭! �tΒX]��y�g����?�S$|���D�&Y�a�#�c�Cd{��SO��]U]�"r�Qy�o�3km��L�(�T�����yHT�b�58:>��y�����ʟ[g?FM��#XI���N�ݻP� ��L��z(A��ⷨ��l6�����5Ҳ,�V%������F;�H]�I%I"��F���FO__X�̖��2�}�1Ǖw�R��!���U)�jlĔ(=�
�6���W�mH���W��m��>���6hҿr?�LO�,��U(,eE�v��$*i][���.����#��[�$�d��H��=|� ժHH@"Cag���L{x��`e��PWu�N2�w���C���l�N�/$ML���F��)ۿ�.�\XWƦ�h=�1jD�X��~�'����$UMV���M�3%��KV\���n��s�.\�$/Lg(隘�P#��֭���M9Q�%]]B�ߋǅ�W�MtiI��צX�Zt+���Q)Vs��P�ڌ�l�e�F�(���L��f�����Iq-#aU�=ϱM�Uw��	��˕]]]�9O<.�2� ��shh���1��߿����c�a
�t)S���{̼6+���7���?�+����Tf�Y�=��Q�7�;mr"x��]"�z�/R�{M Ғw@'d��Me�)��Iy��-��V#Gخ3�:^��FaI����'	�з\/.��$ �@���矁c���Y�Dh���y4vi ��WR�_�%A����������řd�J��$��ŷY��ᩓ����85�w�/\�HR�@3���F�@N�X]P]�U��a@��أ��6��L\Վz��H�Ȣ�^ Cah{��/�4��v�o�=b�U~�8�V}��ܺc�!a�>ޚ4Ҥ�q�Нպ�� r�����ŕ���ג&�w��!�@���l���wAh��Vy�����e ���{	�E�L��
 U^?���Oj���e���d^��X!Y���A>�����U���l�wbXe���ie�;�;ߝ6G��-"�D���t��m\5#TG��tK�s ��^�����.?^{����E�'��/�^_g�Ʊ��7���:�1Ҝ{d_g�6���� �تb��n��aX�l��wե�7ldgѷ�[:���_�l����:�?˸�T�q��Fo��*;)�dWݾ��ۗ�	�����r�Bu}���jĖ\w���,��<��V�&I��g���޾��K)�j��[ː{�f)���G#o�Q�[*Khn�SF��bSƐE��7�{u���/���5�{��I���p};*(]pWKKK3C���H�W~󓒒�4WK"\�Ao ��&�.��`�y�͖�_��p2����^���>�
x_����k��:{���,�UI�ծK�Z!&j7l*JE�!��{Lk�F��eKh�UY&|5�1SV6?Y!��JrM̈���ϨԞO����z�q��9���~�s����>��m;i5m�b�����<��1V:8xb�7��v�tjM����D��֬:OIi�>EԸ�:��'���� ��C/	�xY�@狈��q���|�l������`�O�i\- ��a��VV��"�X~_���U<��ժx�ꕺa�%�5_�Y�nt���P-�i�� �����m�<��Z9vԄ����V�ʎ���#љ`ܿm���ɓK����|���Z�"IDdB�k��RV  Q��V(;�=��?N#�F����3�P�:���Q�]�����%U&-ak����[����*�&k�e�:������Ky�G�2������垵>�˲ϪV��͛J��Uك�K�\�>oOBg������,c���a������|��R���W}0�zo=�R��*�b���9^������}�6ZXo�	sss}�OTI�g���6zߙ�d��������?���Ʀ���ޟE�,���0�`��q���� Ͻ:�'E
ceX� �N����W��Y#r;�#;weddp���Xu|�u$8D�oe�w�t^k���񑊢p�4��Ȍr��v��ך���<[��4F����}!��C�o�R�����ҜY���$��)/Yb�Q;�q�d�M憠7��LK�`�W��C��?h���u���x�N���p $8��d{c���CT{;��� vˋ�����ԷZt�����|aAA7�Yw�j=�����^���G�\�w	~���?<��0��9EE�ny�%�o9-X�^��"WG4j~�.��aX1�$���w�lF�լRF��S��̉�sUw`o�<���:����c����WR 	�ʞe���3]N��'��3$��֦ӷ�c@t��I1��8�&|T�33�uLL����9�->br�ೌDO��2o��8��a�����D�w�*��T�ZB塶��0L~x��[M�y��DNU�ji����0Ps�gRjǽ��̤�����224���@u����b�w�Ђ�z4)tJ�����7r���_�<Hĥ7T�+
o�ҽAu�e��ޱ�n�n�̺Hg&�t��gC3ק �m�JUz�P�$��s�����^3d=sV�i�<�����O�j�Ε�P��:���`��W]�h���m �^q5�jRtEK&l��^?�SH-.�t�i��6K�dA��O�3�dK�C���,�G	h�o=t�d��l:�:��G)~'s���w��a������߆\Ď����&�g]{-����@��[�ze����<K
��[�0<��	h��;Y6+�rk�N��`7�|�t5
���ދ��-kҺ�KG�V8��)����|P=III�+�B�OeEuR�� �BQ�F�͜���R��ހ6�m�2j�j'�<Q�娶,gV�Ը/�5*F���GV׍����K
mnM��&���}����.�v��{�(� ��O�2����Vy����,��P�*�7�������p��R��͒�N�NN�u�M���1@���0Q��8�s��ɲ��yj� Z�q�I��r�A����}��c��T'.��H3"��v����#,r��lU���_�x���-j�0�I^B9"�qϯp	�Y���^��W`�U�,m'�Cy��?k�ջ�x����3�q����(�1�f�SU[	UIL���"��~S��P���YR&�|�ƍa{���`�u����,l�џXmJg��Sp�\+����*I��IڒP*./�P�=z4��"
���$=Q�5��}����E�ў��D�s_��ʴ�Աaݙ&T��Ú�e=�>19�Z����ʳJ5�cz���k4#�ٛ7k����}�@/�^m�����3�X�b��Oa�Cp[�o�{瘟��~��z�x�Rt�\�W�ռ�������[Bb��ZS�Jۖ��|�,�'� ��"�z��O�$��s0�OPE�N���L6&��W�A�l=�yr�c�T�I��YL����p騶��	��=��H���y5��\��J�k���є�w���8����m2c�!�(�G$��f2�RMM������߸��h�ܟ� J~I8w:���"���}Tue��A)�ut�^+E��bܨ��ة�Ey��.ac����q�/���Xl���ʧu2#�������i��}���$��bά��ɜO���!��ِ
��m��%��o�v=�Ǖ��:�v�k<"Fth(���7���D'�ʕ�#��nPPV��O�=j� �t��3z8�3�LI{*�F"��$o��*g�Yw������MH�^~'�֙�Lq!���AZ���yů�q��F���[#����%@9�� ��>	;GiկE-�~#� �26S-�Ru'��������5�1N��;����P���#=^�fL�q%5��Q�|{D4Pb�~ۂ`���
����s�����/���WX�u|���Z���&a���Q:R���� �zܵr�	V������yZ�E�L
3
���E��}XMV1e�2�)"��G	/�i���UUU-+3�!X��ږ���.3@��=U�B�WWʎ���~��*������9/�6�w�X'�#��~?�����Ě�~�5uW��0�t<���i�Ģ�����V����AA�\�hRT��8r��l2�~x��&a��sHb�Rx%��3�����e�=	�C5 =�>�m�I�D+K�;R�����j�lf�q`�)����pR���*�))c]H��R�֯�~�;;;�w�&�$�~�r����i<y�4z���+�ɥ��$�qz��)ce���<y
�%���S��jN[,�rb���e�|�Yp��#
Q��y�!�E�CP0,���^�!�+D��0�}m�a�42�w\WiZ�"�>��������(���ݯ����whq��}*�j��4z@��t$$D�?������{ /E3�r������7�P8Lp�_#B��H��-=86���<��1�
��5�f����
�t����4��?��85;�㫼���������Qi��\��I$��?��]]���.U:��*�l���.(ժ 
/ˋ�%���.��. ��)t�s�:rҚx��Q���U�_����;�w����^Ƹ62�����$��4�L����D����R�쳈����:V����$"��Ϲɔ�F��	xĵ��ۥ�n6T��w���f5��H�(�(`�-*�]�k�h��s��P�Coh����2�S\KX�W���9���;Od�t#�J�U�����Ƽ���9پ��	�K�<inJVTpf�'p�)|*#|�Wx��')�K��h�U��4|�<v��/�8��0�`���~F1���!�6��GVX�🩢����0���*ݾ�bRƻgWNbg��!�s�<�4E���ٳe$ȃhJ�9�!Ϥ*�'@i�ކ-8�&�6z?��A�w;��83�ƪ���B9=�":��p�s�Q6	�����/G�ߕiU8/�x���J���xCr���l
��yoE[4��[�S�OQ�H"ﰋ*]�Gm�6]��IAl�|{d��c[�0!��^������222���������+�ܷ�A���]��4O�a��ĸ�&���i��U>W�N$ާiwϋ�W\B�<��H�H}�<	��{�"��'˚��jG������:�xI�3{���v�Bx@9���硤ÐF�[�R�Z�����
��5V�qʲ�J���4gAC�#���e�7�m�ڷp߃U�8��T|=nlME�-x���n
�b��醠��uAT8�#�.t��E�Z��k
We�F)GU��2�;����pU��	�fdd�k0*ðЎ����D�08xb��%_wfrމ:�q�(��E�+^��F���V!�I.T�LC�<�D�(.Ar�R�#��̆*[+�D<�C4�!;0���_=�,|�|oP}�hX����7������������_C��w��1g߁���y�V}p٩[��=n�se4��%J�q���bצki�6S_z�����[�C�g�����+'���3�)"��W�R8D[O�$�i�C��H>�	z� �ڦP@^��r��\��N�~��+ܙY7e�˝��� �}�bPe��%�i��C�K�1��]|����pM�y�Iq'�!������F�%4��^X}Q2>�M�|�A���:�� ��D�
 ��w�����<3
��'Yr}���v�N���.!���X�kA���6~{��G�_��0�R�V�!�v&���4	 �b"M��"F(s�)�;���~d���Ǣ˶��P��<Ve�Ԃ��U�6N-��,���,B%1�J�<\+X�y&�Ə$XG�}�xѯ�0c��5���ӆ��՚F�=t5��q�%�+<�#�!�B*�����Ţh��O��d��.�+'tkjO��w�} �A�B����8t���}e_����(%�S��m}Sgb�GQ�S����t�G�W��	�`�a�̢�(�O�wSl��pf�踇V�6����[iuGx��c��F
/:~j����
�����D>��d�yH0S!��\�?NA�Co�����K���eee�2���n�e�����T�U7D O��P�o���T��m5����uL��z,"L(�&�	A
b�o՝%���ҷg��>�✖�b�F�m_0�)
��n9{7�t'�/:::<XM�>9������#	����m�7��'�6��F�x:(����	w՝O�v��V=u���Ҋ�	1����]���bi�"I`����=�[b�ne���}U��h]�w����������{�x�^k�uf�o�i�&O��a�D��@�'�'�Ξ����?b:;;��:3��RTkFm)i*e���9��DP����>э�RS�,������-n���7��Ù2��Q�,����I';��4�+�\ƺ�ƞ[���S�γ�;T�b<�4���>�<}�Y/�ġ��S�)ൂwF�C葬�Z.���:��`�)FN��N�9� ލ{���S?Q������Þ�*��2@LX�:�K�؈��������U����0 xI����矑i�9X��r����r���zo��U��#���
p�5>,f��H�aO�U��Gp����F�{��xD�oe;3�YM����*}�W�jb�C�����>����cC�%�ư.��tnE��u����Dk�\P����E�f��r�R��𐀁�>��3�������26���ɲ�|��ѣeD6��^NX��`�È�)���85V>��mË"ݘQv���;
���!��uҀ_�j�n��u�Rguj�t�:����݋�9�V�K/�Ur��o`�=%A�*I��}x&.���:HeA&��z�3%�mӸ�(j��&c�㙘4t�B:�����%���b�~��4w�߸���ۼ�ח+�����jb�f��KJ��1o��0���YUM�%�R�ƛ��k\dH�bSVV��f�?z��DT;6QM�୷F%��q�9
�ke]δK��Jk�=�A�B�:^1J��3'�%����;�'����jjjQ�������ZGVy�Փ!S��a�X):�[�r_ J��B��`2X�<T!��6�'�^8����m�[+�2��buH�	�d2P�Rإt���O坡p�.��S� 9�r�N͆x��݃^%���)��x��؀(�<S�hrRz�귭 ���((l�T(��fCp9pq���M�
�Jnz���
�_bhd�*
�����Y���S� ��:c��GU���xQ3q3������rZ@!'I�9 	;�ѱY0��)9�����VD�Z
E4��-Z;�Ŭ=3����Mٌ��c�g=�(S�i�ȃ���3�3�[t5%���P#|�P�S�D���O�������&�	YQ�{�c��O�&��U��C�+��	[�%;��Z��\�MZ;�"�.O<��r$E).�B�TS�q�Y��β�uD�~*��QV�q
�j� �k&����Ϊ�4�O#�mr� �,��*Pt20ټ�'��eH�2jϒ4�ݙ���E5Y"����H_��W��{�NٗxgĠB0�?HP����}"�B����Î#�zI7r'(�����w��K�o�+G���/ڇ��8dzOԖL�[9YN�/��p[��EeEM���2F�����Y �]i*�9$�i�5ˬ��pz���]��̞�6����ǲ ����B����A����U�'߽ՙ�P�w�e8��h�F%\�����`���7������>5�N̟�D֟�;�{�C݃S��ͪ�0��:�3k��C'�y�Z�L� �nKE�I�PO��
���ܤ���GqK�������A�ӡX���8t�it����(�y�:�Y�[�N<�*C㭁���D����	 J^���_ՑU�9x��H`9X6����ה��g�������Z|d���qŅl�sfi�Rܕx�F�����09�>hH[���G/齴V�׼1=���� �tr��diَ���)n�įK����������baȢ�2h����8wG�T���޸�s�9�O���^ e&�Ō��vD�t˷/���s��~��{�/��?߷z�4����1~MR%:  ChJ'�״:�iܘ��J�a�������ᥓ~|~x����,�*ײ2OkĚ�6�z�&�=�%7��Wŋ���~!�>�=��h���l'd�HQg�� � ~k-F3��M���y�vy5	g�v#�),�ܝ��Qa�$(�*거�*lr��EQc=J?��֒����2�E$���3ڬ�#V�d̆�J�:.� QT�f�r���Z���9��N��K���C����j2{�>�y{�F:���� �Q�G��O.�iʹ� A���O�=?��ZD��o�^&_�������d{�IԢUa��y&�������a;���ܫ5��-�aǁ	QQ<�Qd-ՔM����V���`}|L̤���s�fY��s��2��99D3�_l8�����ŷ?��;�_X�>d���ϬӴ��b�N>	����<ܦ�'Q�M�xPA3�"��,5�=��>u_D1�m%��x+^X�4�Jy.�!���@�l�`�Qfi9e��a+	�lk�]�!�\��
�}�/�FN���^��D$��x$�/�`�ݹ���Lï��/�<�z�)�l� ŵ�b����amw�n�����e�\�Ԟ$ʕ�^�<�`ERhWޘ�����S����f��1se�&[X{i����a@�n+� �O��qi$��>T��y�(�C��?8����� Z:�|��ŕ~�.YS姇Ԭ�"iM� m�keN��������ܫS�r�H�� ;��'9��}�w�P����f;�@ $���y)�CE%�5�S}�&1a���0��C�%x��/�\s9������н���~4��C��d�3�O��%�B�3���[݄
�O��s�;F�OQ������Qs����vN�% ��}l>D��Y���N���#�	�6>��gZ[�Eź~e}��`�Yu���n��7x)^A�_]d�SrS�о��Z0 �K�9���%ɏ�Ŧ!'�\�}����g;�xA��4����&��a�Á�!K�� � �|%%�!0�[F�S"�umH�6V�=�-�l���Ҷe�"MQǒ����׾ӈ�_�6�]��y��t>���&-�����\I5��L͗ˎ�O؝�{H���|l�sEU㐂D��2�����T�	���n�)�s�K:n5=|�5�j�
�S�d9m��������;���_.��]��(zI�l�@ x�툰�%S�)�1�[WI|�>�����M�c�	
R�4�TKu�š�-]��mn�&JAոY�(�/j}�Hm��|�����d#�l���VS��rc¡)�3��1"�j��;/���QE�G+zo�;�祩��hz�Sz�æN�3%�a
��W<L���D�1vr��oa���`�J�c�	�ҧf����1�I�<�v�o����z�J=��߮g'�)��^Y�g��z��=����L>��ٺ��|��Wi�����e�=�h�{g�6m�g��S�mT6�1���b�����[�,� ��zE���ٗ�k�ƍ�+��:0�^^4��M�y�����KMY�����s�T��pL�pƚ�U��BT��|�%�ąr�zI���}}��ϡN5r����� v��%��s�s:ЃBq��ь�8n���t3gcC�w��é���
{�lv�A��!��:9����$�Z�e�XNrr��L ��U9ˤM��Q����٢��^m��-Ə�Wmnl\I���:��,϶�����_V��5Oϸr��s@ONY��ng��4������R�����`p]�z �9�=������;��W������l��z����%�v	n9l��+���0j��H�P_�ߦcK��ը?�xÊ
��:qbʟ^wU#PTuwBX��<ĉ:�T�������5�[b��t(���o�ֻ�:M`4>��mhhh?�]1�4�n�)W��<��?	�b7uWo:�U\A�S���[G��DG�q-���ׁ�h�m�*�#�1�`�3�5Ż2���3j�Gd��ܹs�Z�'jgN��죫d�_�r��N�+'��%**������h�i�]�|yM;W|0�H	��E��RoUN��e5휰*�b^cO�_�p,Ɨ�򤒶}��td����H��ˑ���j��z����L<Cƃ�R�gg�n}� :*��|�W;�BM���?|�N��W�u�¿ ��9��]$��¬��zc`V
�ޥm6�D@��l6�X,VZ��t�=k��
������~�E`���sl������kkѥs0�Q����@F�[1q�����3R˿�Wڢ�{k���h	�->�*}�]����:xt���J���С9���"���,֘��@��㬁����Tx8��0�rw��x�5��^�2)�<�Z��t�㜶�mAq��;�R�O|����U\#��O/.h^Y�nM�"(�.`��Q�С;W_������*`Z���Yf��spp���Gٚ��]m���,�a�0�g���G����E��ҋ@`�z��SyrE��)}~�U���zm�3]�Le�[|�ӭg0Nh�w��	����|��N����=_�N�$�t�\Ț�����������掵��E�|�v���l�b�Z���9~|��-�>���1q�9 �w�D��K>����׾ը��[���7E��t��56.�F�=�k�S���W��i�:�/��֫������=��:ڃ�TVU5o<���݁��?��Ia�qo�<k����_�~���:T͂41H�������*�.Y �����jʜ�oI�I��]���1��o�3�J�a��U��,-g&�Ĩ��+��w�|Z��|���55;�"J��AS��_�+�`�kq��+���|)�M�+.�	ɫ���6�`{u�������mU�;�.�F�a׻7�Q�7�V�0++�#��r��LN)���}���s�!""b�����yn	�������`�N}���7���E6�Y�l&�������5A	_��h�?z/���{DŇ��P���} ��#��
G�m����:�a?WX[�<�b�Q{���h�Q�1�|��o^V&�J��S��9�aPĉ�+d�,������5"�ɏk��r�w�����9nX���]VC#bi��ׇ�֑������q��h�����4G����|����X��x��tT$�}�b��Y�T��#U�{��3����O|Ӆ���jEM`N� �l3��}[C�L�g��O�x��(�]j~iOfݫ�999�	��V	���z�f�6����9�VU>� ��\��V���V��^����jL0���*������-�+��QC@�W�,�F ?�P�?��s�t�����PE����j�Y���z�Q x��\��Y�z0I߷x6�Q�R������/c(#��~��[�n_�d��9��4ߪ��Hڨ����iG'��(%뻎_��)�d��!���o�Jl��O���&�<T�����eX�L��7`���f���rT3�{��"«�u���x,�l^������� eʳe�+n-�S�}&lo� �.��H���������;�M$Elfqs�B:�DpO�u��+an�7Ŭ�ܭ�dd�	�4v�Bj3Ğ�Z|�!>w�'4)���}G����x5V��L�E�=juHc�}��`���T`N�S�]�W�9���*���� �J�k��ް�c_U�v���] ���=���M.:��|����>���7>��0�D|�.�����〭�]9�
����&��s���\d�!�6�C=(��x�?f�e�?�k���u�_�;�Z[++q'{� d��v��xy��ϲA����J���Vb��J�kj�m�D�(٣q�t͇��̔A���E9�	n0^P�>$�= O�_���U�K?�k��a��Z�i��,bjr��$U^��b�NM��N522
[O[��>&��ba�$�gL����^�d�*T��t�Q��,�U箜�5S�Ź5N���������$0�zW�x\A4�_��+Ŗ�Q�^����n�eB�'�{��9��a֧v�^�a���vĚ�~�L�쪇J10�߸k�ׁ��!�O(���p��T��TΛ�L�qzʼ�PCXD-��!#�n�яk_��:7΂��ǆⲏ��3_	�{=�)<݄`�G��7ƾ�kX�a�4� �2e�e�����O��š�:�d����<��5+���������W�C3FEM�0�W�ဣ5>.=NP���"���ُ>c���C��9�->��!-!��h"�0/O�
^u)~��y�Eb�8@����%� �ѕ*�E�/h90���F����8l�[]Ǖ ���ky����Y�\��U��fi�XM��w*�C�S��[�5=A�)�k������ǎ}��[��sE�ј,a,����a�I�w��c�޿��B�UT��%Z&�\<�u+����'$�^to�	9��y�.m�e�S�'g�[[D��4u:���Tx곝>���B�c�����9���m�ҎJD��!�����-�зʷ��C�������?�2��K���5�L���Rw.8twk�Ą~F_���oa��Ă�g2&¶�_��JT�ާkq�0D��v�Rؓ����,B4�|C@�	��Z������n�y"��� Kz��>�E���̧ͨ5� ��?����^Q7P})DD�7;��͖OT���[�#m@*z�[$���^�g�a��!�N�[�x6���|��V��h�m<�@�9
e@���J��].T�w$���������/{��@�e���S�4@�7k<h��~jR��� Q�n�Z��d/��gq���;G��}���E��F� �>��l���f�(� �WCv`<>\��ϣ���_�p�R��I�xڴ�n|T�_��8~H"�d����nfY�XO��O���L��)�Ji!���r�3�W�9=��E���ZujKcc�����Y����ѿ��A>�\Ƹ�����B�l�<)G��if]$��yc�!�a�$�wN����h��:b?�����b%�o������#�[G� Їu�����i����E� [/�>�����_�R�c��N��n�Af؆�V�ҝ �=���k|7۟yFɖ�T0H�"Wa0�m$E�p4�80�Y�G�"�e��Θ�g�u�q�������Y�Zpx@�yO�NC�"��;��3��w��\�k�dpd��*�����gY���2�0Z�����|�V��(j��'�jh1��P$�H��ݫ���Q���c= ��@I7�+O�--�]}����S/f)s�5�a����s��
AWP�m�?����X$TA�&!^�0��ڂs"�=|4��v�lE��5��c�2��7:e���e >C��k�:^g2*�OtD�&� %$��>�;����A�K>,�c�l�t�mO��?��sM�/�,2|k�����b![�3a����W��-5T�o&�p@A����B���'A�-��yF%���<$0[���ij�$��w�2�y�Yc��C��\y�/?u=����Z����"�V|�]���M	�oE�ſ�654����֟_�5�{4��|Z��b��Xa�������X���A�7ε�<d���*٨��,6w��z< `����SBpw�m�ft�㢅;�f��/4B�1��{��Z�ۢ'3[�f�*s ������DX:b��uv�R�g��O����=8PV����$�G����$o��\��;�˭���#��� m��3��'�ː�?�<�j��~x|�P�<��?f*����߽�@�a���_SSS����UU�Bc��Sp^I�����\�e����g߃�Ao���H�
�gn�p��ݽS?�S!6��>O�Վ$�6��Q~�R3�m�E�/�OK�: %��"t��c�e7�,���u��sy?GN=�����f�;TK�sE�
>ɰζ�v<�:����hs�������� ėυ�KKK#���5���n�Sqїa�-�{@���'��.{j�Qyn�. ���N}��Tf����8����R���T6�6���lrr2�S>���	�	Hzh�P�wۙ�KY�4n�zd�ߧ��2��㞵��Q�+'g6:��O��4��$6w�yn�qXxVUn�ӧ���()7�O�ސWC�Mm@C�Ω����oU��7�K-���s��'���rq�6�9q^���������8����(7�c��ok�߶�Ց��X��b��M?�J��a�gay�v��w��֏�}�{ʭ���^wrx�7��Ƭ��(//��D�G_���dJqk��h�&�I>K�V���a����mf����r
�%��N$��(��	���S�kS6/�4,�3��-J�홥#�������;�U;����?�onf�G�U���=m��7��[�u6�/���*bU5�����S�ڈ|���O1��3�����ò�k/���r�����»��.A����34+��އ�u�^an�M��--��K4�9�}�����ˇ#1ކ�ĞY��|��6�K�D!	�턌j<�"���(��`X���m2�ֈC4��Ի~o�n������%r�r���W����u�̡��:3��ݶ��꠱�����p8�v.�s�F��%O� q,)j�N��pG-at4�@���:�u�=�wvm��&//�3�����x�_ uL07}|gz�u�ŋ6l ��2ɣ�(��sA�yZ� uŚ���%T��oݛe��"�D�z�ԫx�W �����?����V�&
b\�S�x�[[��瀮{`M �\o
'��oߍ�f=�Ռ�9�p����L`�>S�bl��c��F��ic~S�D��q�E�od�]��'Q1#�+��O�eF�RItf*m �����x�C7��KZ���*Ugg'�e�����ғ�{��Y`;1{-�)UҾ��;�E~�KPU�����Ղ��6`��#�b@O}�=@�G��ݼ;s���O��i��|>}.����w���ā�W�l@�O��{����^��A�ЎpcQ&z/��K�-�_����Y�(J�+	�6Xj�����f%���i���ɔ'���B_��aԪѷte�V��f�@�LIsV�Kq�/��&wO:Y�i%?=�Efe�q۴v���(��6�\ǒ�#&�J�,+E�Q$��B�����۷��X��,$a��k��}�Ѻ}�a�}��n��拣�.>�Q��26
��oR5�XtS��Gh�M7���5�XJ.$�#pD�E}���{��b����Sx�"��fѪM�/�+V�-¿U\��B��!���g4�L�=��\m�筌��HBK�`��/U���&S���)�Y��x̅,�����n"��v���Pj��|�����R�鋮~���?4����RmY�g��.Sr�%���������,nCۊ�tޫ�Ј���b��F$=/LLbs���L@E�{��% ��.�bH�5�F����^@q >�$����©��%}��j���-���Xb���>7�3מ��OoJ�.��Z�|�ՆsV�Y0�����8}�׸��������z3�_p�z�� ��C���V�1Vn�(}�h˕���:�|t�y�Hש�HVTG�*�.k�|�����y �r��0����o+i�m��#a������r`�R��i����+`3�@�qXwWmF�h���zgK��;�Ô�[�����{$3ِ���z~SR�ˋi5�
a:���xj���%�ag��D�&L��>���o���o����D��״��#߾���#
2��]���aO�Ё�Î#�w��iU\#�L�W -��-��ۮC��V9�e�3j[�2}"��t]��j�si6L���׼�
3^IM5o\��D��D�=�'<X��������?=�cm��|<�4*��D�����5�0ֵ�����4L/I��*�4#[F��0P+%z��*��2���5K�W9z�5�����Ukn>ѭ{���Hߒ�鋸�6`;vR��$W�]�4$_3]�q�E���f �>�5^Ϸb*�y	��*B賷��\r�7Ӧ�=�Og	���oq��px�ӣ%���/��������K�ć��(ˏ����Yk��?�9[f��&"��o��O?��`�{�B�!�d�s*li]�\k��6�h� �?Xg�[��X���2��;��Sɽm��<����ʨqV#�$�#�d��jj9�.��Ԫ� X�	��Xj����������nA���S��E�da��|D	�F�c�0.��nq�ʕ͍���Zv��~R%+6&� ��kl�f�2�m��2��eM�Ϝ&Iv�w��-��󛖎�5���-1���y�w��j���׫�-�%.� O�O���H�^R�LL��h,���g�w/�-Ci��˕'�i_�~�n(xtQ-l�|;�����vʪ����$&���40TSS��� o�����֪���\d��羰�(�K`�]���܉���i��쨝�3$�I�JЧ�9��� 3�E����;�������^3��\�w��'gQ��%Y��>؇��ދO�=�Pm���%=݀���(�J���!�w�b �����e覱��;)le޺�N�Q���i�b^��#�W�9��cS�E��b�a���?������i �\�:��G~�1�J�9�o�32�U�Qt����cR���L%����hƣ��z֖�Hp��i{Z���4ι�$?̐.
hD6�H^c�ȫWЪ�ޢhsӗ�z��/JQ?	d=`�K���ma V	�$�����?�޷I��뷊6P��
�@�n�"z^�t��M\ۥ��[P8P�o�ð�&�]ƅ�K�j���}�E%𫱩����D�VVi=��i��'R�[5����i�o~��n���3m���\i*��}nS[[��}��-�M4M
Ͻ���D�(��˻5u����$�~���	�l�Ot�@� 2��*�0�_ec��.O�}���u�*�챪��_/���a���i���%WA�f|�{
-p��?x�����������4�R��=�J1�o]�^�e�PG~�iE�]V��^'��h�@@��<O�[/�������mgN���zI�=ŏs����E~��%�&����s	[GwYtU��e`�Ex3^�'m���u4ʷ�Bڸ3�z���jVߠ�;�#Q�n��r�.%]Bxs�J�o����|?_�D�����ی����2�t�,�L��*G�X����`s�;��k|l�Ľ@����� @V�RAmLll�D݉��sP��_���Ve���/�C��^K0/
Bꨝ�I*v�FAu�Y����WH��8���-舵wk�\DI�16�r�s��G�����k�d����X�qȸX8n��6�_0�?�j���*�o�f�����N������6�G�����1v�r�>j[��vO�{�梧����&�!�ֆ�}yi5�U����f]�z�@�P��I���R��ʡ+dź�uO��[���̷hdEu*��q�K�����0�/��mz;k��C~N��c=�͋=�RgwW�<�3����o^z�OW)M8����9��	m����%���K���a�s�l��ʂX`/��'�>u��ǟ�jloqȉ�	���I��]�7���8�o_��^��;��Li{$����rWa�;���
]�ғdQ�Ԥ��д���s�K�r�f�t'��aA'yYS�g�M:�k�Ӫ[��#�ZJf�a���/�{׀8��b���VG& 5��4����.�'N�ߚz��:!q��OJQ�ͮYkvѨ!�H�xZ,�������g40�F#-�#w4湣lv��^���;m>zD$U�/QH��l����QHi�����\�v	'��^H���~�e�Ι������R�� N��	�~̈́����^�ky�M2���qzv	bV����掠��^k$h��Ol����6 D�?�S��/�����M��Ƴ(ӬΗ�C��d *�3[tX.t�i�z��Qlу}����e��&��I�89���J)��� ��A�V	l1��y��Y6=�y-��H�f��S��!�ʳ�gX�,���J�� ��tl�Z��~�����Q�������G�a�z�9��$Q��6?)��ٷ���v�3��e��'����t���G��,�P�6�؏�7!���G���<7�W/)�k��e�D1�#�F�|Vp�i�}Ǖ��U��+�P��!��~2Wô���͗=ܺ�Aݴ__ML���> ��n��џ�+���g�>��m[Ŧ�Z7�{.�<�L��T�W
�T%�����6I:�|��*���!f�u���@�X���Ȭ�T1	E�qK�*��[��4S��FcKJJ������D��<��b=�ʾ��^ZY{���$VT��CM�ړ7��okU�&�d�~���D�EJ�{�Y��J,��T��G�����4&��	�f���7������Ж|�5�V��vѹd���r�Q�$����i->a���њ�c��%y=.�����^?�"������Ӫ��
ccb���g�iX7���^�;��TZ���ya��ˉ���L��S�GzY�0)w�z���s�Ϟw��L��}9xOz1=�UP�X��a�J�*�Y�Z���pA=ٿ�|��އ���o~a�d�4�Q2y��ML�~8�݂=	��>���WE�Y�\���� 3��eѪ;�?_�X#����
��DG�Ri���j�؇ر{�����^����葱-������{ѫ���3@7��`dd�"I`�9����D�~g��ק����,����z��0n��&����r�h&k �����1�{�Z�B`/�e$��;Q؂���-��W:}�6�����r�a�|.I�a����A�BOks�XE�uD�g���&w�	�l�ii�-_Z����5�;��x~�W��[e�6x��<��u��Z����8��,�@��}
$�$�5iHmmmń�u�r1�Ʊu���.��w ��So=����h�ތB{��}*o�0v@Z��I�A����H��j�k�:U>vw)��9f�����R	�]8����M�B�/9�T
/�u���_6rv��11����zI��#dkc��P�+f0*��L�־E����g7�M�
�$oF���d�������_�X+eM%ׯ?[[[{�Y�l��$ǝx����77��n�!�ntZ���9������> �[��/�.>����=U=��ө���a�q�U�?��v��-�߆�<���D3`����Ci??�;�7z��'�хz�y�&�8�ۡ��i���̺�VN�x��O�e7N���G�;ɖ�� Qa����řu��U�CPM����x�.�
�Y����ɦ"�M������ �>�^;�r���������L���
Q�IyT��{���-���$�p�N��T)�քƖ��#���<q����jE�ŪJ�d5�X��.O���i���C���^�9{�:n�r�=Sk�@�9���	ۿ���(��J"��Re����2��j٤��u��n΀0�"��ҳ�3��袍����J��lH+GA8���N&C�ǜ���|����C���I�Ɲ�`˅�#�J'٢d>Wa�K�Q��ѣs222ȧ�Q�������]X�o�V�B^rVX��+=-�{X %�h�[�<k� ���Kh;�gּ��~cz� ���Z���zzz�aއ��X-Y�d�r;t���O�'L?�[��*-�߁~��F�o����$"�=��ڮ�(�?��pF'�,���A�)���-����d�b[�Y�z�ft7�"2z�sŖ>���m��3C�"w"�`��#��Pď�+�D�������q�ϟ�*��0Y[?[4���v�`4���� ��*����3A��y���{la�aa&���c{���q`+�������He�:��!�1��ϣ�Su���Qm��Y��|���_���{->���0�0m�g}��l�W��nPį���z�9��x�+�AN)r��K�zѦ�Z[ցj)
����]����E�����"Ǯ��Vw���X�}a�b���2~���?4E�u\����Dk>�]����$*��;d� �MV��X��r�����(
H����Q�s�-��mH<g��BZ�c]t���}˚#���B���9y_�
�	t���s�-n��ϨȬ�CV���B$���s'[K�N$V)��z])���fI�[������7��Jŭ�F��At��H'���&�N�+j|���B�E�������%---L9�k���f��'
E'+�
��� �������������gV����$yS�N�a�#�Ƥ��ӳ���S��#"u����(����x�*��������;e8d|xd�ī-3��Z�#l#���A���2Tў��
5�;�h������P��]�-�~x�B���p�4�Y�����59%����Yd6:v?\�Ԧ�3�o�o�
������R �����4��'걷����B)Ԣ�'��_�8��� �rE���<
S>��8�P��d(�xEQX�k���ˎ8��l��ɖ˫7ru���UU�P��$U���Q�OS!�mȮo6�E��z�.(]Џb�d�(�!�������<�|͉�Ԣ��������P�j�3�EY�K�2--���N�]EGo�&�0��s��@]���C���)����uV�*��碉/`'�NVh� {l_XQ�u������Kdt��G��xg;;4S�&J7P��W��HI1�te���/Тqˌr��\܂J7���i�!<w�5~�8�ñ
��1�B�;DKW]%�j�Q�Nܧ̳���7e���y�jVU�H��F���)�K�(O>������+m�O�,��� |��xqޑg������@t��	Ϭ@��x��*�����m4�-��l�
]~���'�?x�G�?kl���f"���u~�z������Y:�fi�hB���46����4��Ю��pg�a�����G/-���$�;�`(~�%�G�G��y��.���YM$���ڬx������XX(����7G�@����	���i\�/�:0�?V�wt�CgW����\�O&:w��B�5A��m�����r�$����F�j���.�e�C����Z�S���)
�i�����L�|Lk[՗>0�_���#�s���$��>�ȫ,u(O3��Dߙ�K�s����-�{�LE�5C���F��?$hžH��	"<���n�ZtT=�iH��16��?#�Sr�����Q.������������݇y7�Hй��V���m��-Ϝ�b��lї��ʭ��P��?��-��Y�~������|��m�����~����$:ŝ��S��-z��.B[x��TbCk/+��!�
t��?VzGlz��?�/B���!�ܤ���O�)Bh!I#�����Y���DY�Gr��؉�����n��Q�u֬v78 @��1`��y+�I�s��Gw�]�]"ww*����1T��D�Za'�� "J�D:��L����Ne���b����l��:Q'���K"�� |�5�5�<���Dim~6�� �����<�ʬ��L_j��1)ӂ�
���74c�THei��.��5�6M%��2e-�a��ʵ�F�O7�|�dO�,ג����������}γ�g	�|/�h`��o��M�+W�C���/���x�+OR�ė�7H�0�0�L��>��7'5f�>1G*]�	�FЃ.#�ơ�i5d�z�p�l<�x9��Z�#a�)�c(�^:�c�7�\�.�P6"+N`�ե����/�K_6�UÉռ���L�/��y�[k�D�ph�_����s�}�4�O�ψ��'!����7}^88�-,F�q��zx/8����CQf/��X�'f�	����э����D�[��s�]��=DF�gp���A��ް�<����T�:;q���L�U�����7�#��7�>�qEx�1��5�G�qN� �+�F�A��w�/�@mvyX-�}!�?�p"��3�|D$�M�0mxF�H�& ۓ4�Gة=#����M���Ygq����U[�>�������E���6�x2=)+n*�����"����5��؏�4�)�>�$�U����c#X0G݅�v5C5��GK9��+@���<J?�=p|��� <�(L��=}�ғ����}i�+��d���t�� �G�Z/}b���,O�`������K^eV�`Obe:�U4�I��?�g�F��Ht�Q����N�;�lobퟯ���j�(dnƱ���q��. ����J�&o� �SMS��ؼ���!�Y��.2��ط��!�/�0�ָ�HI�%��+���<�}�ȴ��A��'���R�Yo��Z���LF��fX�E�Gu�*K&s�E��/�� OC � t.����������"�\'B8q}EQaaS��k�	v<K�p�j�f����s�~�W�����0���a�)�k#�Nk�ʐfkK�-)?�\��{�n��,���2��m�;�����L����]|������4�;���8�yu�Z&�I䯮+�-��rVU�R�>�b�|k��7.��쯠͜�nݺ�Z����ҭ!�B�]��p�'Tomw�a.�D�ĥқ�$�7�ʫ�J/�ry�;I����F#���T��OJN>�*��v���-o��+�R�+cpXc�_��K:�@y�lG{��=������ʆ%3Rz�kmG���K�ѥУ����xR# ً��b�Ìk�VQ����^?o>.�0\t�@��YM����j	AdЅm�n9G����<��$�A'p��=�;r�Vkp_X��Il~���?�c�dvոϹC:����[)��0�:���-��y�d=~NJJz����ZIT���&.{��㘨6&�)�k����?�|�'�b[G��1d�G����δ.P�x`������
��O�pA�)��f}�2ڲ��k��v.n/�SC,01�aq�y	ڕk�XK��f�C��U�� WNM��\Z�#~^l�K��L����Z.wdk��-c�`>9t%��ɝ��Y�Z-�/(:�֑�6}�*C����ɺ�IcўSn���):��*R!��#�a��g��qSa�&�&d��4���� �H]���u=}:g��.��'�-SC�U��.�51�{��<: Ww�����z�MO��M.�W�ӏ���[��~�ޫ�P�DW]�9^l�)yƩU�8���T�%�b&���sԑ���[J�m�G�:����?����_���:�/�ZZ��������L���h#����
<$��N�*./q�}�Aǥ��#k*Y�9���*�W"N=^�ϛ�ىZ�!_���XI���m5�o�"U�`���Ҡ�̑m�ǘ�.��ND>r��ڒ~,�/{���x�2�YE��������X���}V�����=�xH�G�45��\���!��<uj!r^��0=�fO	�	W��i�W
�p�!<KLg�B�A�Yv���Ά���c�Z_�G�r����j!��;�1ٔP��v��s*UI�� �Ջ^~���Ph'.�ҥK�
�t6=���i�!T�u^���!9�z�箷���f7��mz����C���K�ky�HR8�SZ��"6:\<����Y����w͑�!<l͟����655��Ahr��}�����Ͽ�u�Œ���"�2))�j���)ԡ�e��t�C�kRTEA�h�{S-;Β��_�=i��@7�H��3�����s�~���H<���ɞ����Ύ5��a"�op} 4a��P�����>�����(�1���mXR��$F���9n/Z��[��;��`�Y�^���'� Z*���6�}���$��9��}�G9��V�c̄
��ׯ.& B�_�sd�!�7~�C��rl�1��Ǥdh�.�'9�D(?,����If٨e	x~0i4��o~�|a�L6�\�!�%f�d�ke.�_�Q���psTK�:p�2�z�`��W �c$�i��ƴ� 1�Z���쿕Sy$�vӦMV�h�+T�V�t'@ �z���n3T<}�=[�8��Ra�{�3������o��OGr�݆����⠎
��*�(r�ɉ��-��z���ʰuui/vH����?'��>2�p����QY��v/�{��#�'�)A��[N����=x*x)�_#//��z�϶;:�R��iϞ���$s3B��ؾ�E�I�Atx(�J)�O� �|��@G@��U;�xv��|�(T?�Z*�o1���A$5���)9�9�P���#�jp>Ā��c$�8;OO���p�=n+��ԣv�kU�\���҆&�zAL�å�|}��f�QK�;����h=^�]�4�����Rl��64�9����Y�� N�֝�CI����q3#y�7ǖ54>6�;b�x����7���n����
X`�߈����:�a�iҢ���6�ܥє�o��b�ῈG����F?�_ (BN;�We� �P$oZ	}}�K��p���a��p��L�
n��EFSrXX�����[I�6�=��;$��I�r��S}U���2bwkAz��G��g�c'[v19��b2\dVS�A����15�\��@�+Ɯ̨���4i.�; 	�lG��J�ҢJ��+�����C��Ȍ�ŋ<.C��6F�#�I�����9���<��a�����(� �ǣ�ٟ��=K5w��PQls�w2Ĳ7,	������B���a�轫�pe�,�fN���ִs s�7>�4�"�.�C��Pg9#֦�s��U}_�y�<c��a�H7�i�闑�A��n��XzԐ<�z��)b�)�~�P�>E�t�['�S�&�ȷBrWg����ݽ�raɵJ�F�1�o18\����e��B�bȃ/5��Zi����
d���*�_ �AR�q�O�+���Y'���v-�����e"�P޺��;�M����Zr�E�qN�?KI����}t�{��s6�G�tw��@������4ق���N{��0��I�����-�yO�%�AŸf�?�1�<і��ȧǅl
l��0i�^C6(���}��a��7N�`Q�B91f<�z�}I�etQ�ik����{-"��Ԓ0j�fG���A�^H�!hR���}�hL�6���6{�S�(s3��qWnm�I/�a�NSX��y���E��'܈4!����qs%�q�
:&p!�P�)�¾����yqHL�3�d�E�/�ڰ���&#�(һ��1���\��vڜ��Y�E�'��,�\r����U�u.����E*� �scD4�1��SB.R��Ͼ�����$h��Q;�2Nu���q�#�q�����"1^�h:W���A��I4=�t%2B��9kC��9�r��1=�>ř!3��d�q��n�3J�L%k��C6Ue{_l�GS .�e ���a���噹�X�������͊1]����E�IPl5��o����j�a���3EOq�{fcK/��#M�1��kӔFp��hgV�\�o�@��D436lM��O`1Ѣ~��gVVV���U�tRӁĠ@fn����K|I��B��Ym��ټ��˸�ud�O�:��戠l#�2��o��Uw�����-a����#�c��Z�05g:&���P7eq��"��]���	�Cb� �w=m�U9��Ќ�N_G�n�޿��&�A�+x?�Y'� i����X�(��������xŠ1��œ6[ �<���aVʸpڅ#��~I ��G�B�q���~���|�����y���Qc(s¸���e$Sq)�d�=FqXA'�C	E�M_Q!x��Ny������7r���}k�8�r��"m��9��{�{�v�b���g�2@I���M���*zW��Z_GR��n����q�8�9�/�g��(�!��R���r�*Q��{��������%��lGm�sy��g����F�ˈ~U�🞞Nj�khl�7+1{pZ^G-םC�`���#hH�RZ3�o��J��T�L���w�޹�G�T\Z�8$�����U;g.|�g_�\n���XrL�^��s+%烐|�4ڤ5A��^�%EB�WQ^��.���mHR��� �VNޣ�q�*p.Yg-�⚋�y��Vi=Z�2T^^����&D�o
q�suu��Q7r�0.@�C�fyef�N�+�qaSC�����?!1��f*��2杁g�0r�puͣ4-���L6	�CA�-H[����QXV���}��W�YH��E�)�}��>m}^2$ǔ��� �#H�r�O�S�51��z<脗�D�L=*�_zA�Igd4�|$��OCuS�<�ӡv��¸*��/E�1���﯀�~6�bW-
�<��b@Ѽ�O��?�b�<ŝ�+!rtt4n�7~��]�'��n�%;��b5e�'p��t����v�Z��ND˺��cV��ھq��+��9_x��"#��+Ƿ#�v���MY�¡h�Q������iث��y%��k?,���5b�3G�D�+b�-��8���q5��SЎ/,ҫ:N�,����C���<|՗�znXB�(4�Ab�_1��3���WF��Ν���>�(��LK%��b��lr�6��H����L�H�M����drL'�C��e���f�i�ߛ=��܉�.�V��X�Q}9Va��HG_�u�Mw�{x�]A{A��U߶��$�,:�V�Խ@��1���v\�N�g27B�S܄����vK�E����s�_�i��6y���&R��NU�K�J7����xej�/��S�#yV���s�\��&���gA��k��8�t<��@⫵�Ӝ�L�����JHox�-�����L��3���\���|<u<�A`��C�6Pk������e���'����̼v`͚5Rھ��XF��@J\��6��#Տ��=9�n$�����N�Tˉ��*����&\��X�E��[�y�	Ws�:�~���1�:�ڟ�Vs�(R���&8
t��DA{���o��}�������,֜�|�.v'5����C�?�5�'��{̩ͼ|�ϒ�����4@��M�t]%�3`�R!���/GL8��
n�[L���2)i�S���F��h��w�X3v�;�H5a����Ql��K[T���6p����"�JyX镞�k׮�%%%�29���_u�+�Z��m�뉜��*�+[O�=})�����W�'����Qu�L V���'��O}�^0oNߡ���K������"Z&�Z���x����	�^w��D�փ�DI5�F��ڥ�?3"	l��s�O��HF��D�U
6(�H˼�7�<<<|l۶m���/)s�*���P�Γ���%˶��V��X�8�E!w#X�sI����H/]��"�s��R9Y�CVL;�`m�J9�R�)������A�v	�4��������|nm]���"���R�m�WNi��yFDR+ߵX��z~��Ӵѝ��RPL�籊�v+M���ʳ૘���o_���G��u��`X���ۘS=v�lin�������>N�IQKGr|�a�w`���E?Y:Y����(K�����L"�K	��e�_���+Is6�
6&���_ �:�@��#+B�H���5�H7̙ɲhoǿ�+�� ��~++i"�|08E]E��QY�덷x3���i���)�Q�z�uNW+�I>�{��%�ʱu��^���1�<�N�5�z(RG{3�迅��|
=���qWq'"1r���Ju��l��ҥ��))݇�� 5���qaf��N��5���s�{��� �����_v-�1�6����3����۵v��	q]��<ܡ;�pvv>�o_c1��rP
[�"-^�s��`�%���O�|���u5.'�����zB�F3]����� �	V������N!���?`[_��262�Z���!�;,n8�]���_yj��`b/X�{���Ch��%�����#��C�����v��y�>yO8"DB|i�������=ʠ����Z��}�D=�8��z���;ۇө-�^���,�Ks�b���Ar��q�V� |r��:Y�۽/^�~-w�ĉ��JShe���U�XB)��}��WN��S6,� �A~��~�W'��;l
�VA���u?���_��O�OG�y�0���Ƞ����Zy Zy���hq�e��1��BHv}͉�f��577S�|��nXIZ��4%!�c����*xG��E9L�^�w���6�a��CW���\�KeYݱk�Kw=V��NC~�}�ػѡ�%ee�m�]�D}r����q��V|�x ���*�w��.^���gD2N�Eu�����H��?lN�1��������m�����]�Q]��#���N	�}�k���H��Ojצ����]�a�Id%�D��9�B��hI]|�oA��x���}�ow�)�߁�B
_��ބ
���넿����m$���_������>jdJ�kŋ�05§�o�Ύ���c�l&�	��G@؟�����T���=�D��C�o��߉D�v{��� �{Z��8p�~|�����x���֓�^{�RH�9�)��:��Fڲ|��;m��������ש7Ab%Eo����A!��A*�E��?} ��˸x�@~ժ)�i���d߫��4�
�Z�4|�ꘋ,���WY�Ͻ �Ob�=��Bb��p��Oz;�)���xj�>�=	<l�'t���"�\��r@@m���Py /D��#��S)
�r*�@ĺ�����\+b��^k`�G/X�@�-�n�B=v�v�茋o�aG-���ٹ#�ܹs�UK!�#�([�a�xVo�2�Ѫ�.?��)#"lepFL	�8eK( �TVJ[[[kD�?1�� *�ɾ�n��i^QJX�7r����=���<���cKAr��� %��:�۞)�#�D~[�E��i�s�oT-�x����_��.� [Y���u}��Q��$I�DB�z��&���^��@���
�u����v�lO��7P^2���;M)t�������B	[$��$%'k?x����;���}����θv�ɢ��KH�k�*d��]����YPZ��l�4%�L��Pw�f@^�?���wl�F�B���ew�[G�R���Ű��O͑�N%~��2(�����i�E(�&�����H��
޼W���X���t�L��U'wJ(m��2>:���Ո=M�S7m�!���F�U�V��ȁY�<����L�����j���3�.J�h�� �RGTM�9�W�ʑ������ys��.�h������(��qG��s9�M
Л��>�A?��)��ASd^YS���qc_NUU�-��P/������Sc�iJ�᠂X^��?�OG%��vcO@Zro���c�tݖ�$~���g�hh��\ivе�A���o����pV&�p��x<s�wN�3$X���3�P�!9���L��QwM������\��t��sB�7���o���n3��,;�my�����3M����^��F3�ߖ~{�W�<���+~�1{Az�U��q���pf�dY~�,�?�X5	}��%!ȴ���MSp+��p{�������Ⳑx�z�
ڞ����ҫ��N�Co(�t��m�'}U���Tl`�;����~XL5��{~&�Ͷ%C+�#�P�}z��{z|��)�����h'���G��V�!�%ԲR(��Z��kd��T��(��ʿtW!ic4�4�����y??1�΍;N�H,����d����fd#������)I����7'1n5C�?�c$7�;e5en /��v�^j�e�/B �[�Ͽ������%��+I�/�{���я��c �"�+S�~�)�u��|��-�?Bydi'�6g�$��@��������r�J	�т!o�/���(���YI�4�nN+\�GJ�z2�5mКf5ш��S��[b�Q�?Aӣ���IDA.�6Y���^�wK(��+��f�'!^)J��"K�¦��0��ۨ5bКy�]�6�p�i�P i�]?���{N��)�3��	Y�a?v�œ��1([�Ux �ܼb��'B���{��T�T��d��q�ԏ�߳g�ڼ���Fê�W�sH�'K���|� E4K��
�M��?[�{�L؛�Oo߅	��!���F�(*R}^�۽�nl��ޑ���4h��g��ݹ&1>~^[���^�>o\�7�o�}w�ñ�BJ\�p�2 S?��_�E?���a.Q�v�z�2�6���+�Lص!	w��m�3�M�����PK   ��X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   �sX,�׳A}  7}  /   images/3d46b7b2-3c4d-4bbd-b0e2-e734cbc728a9.png @迉PNG

   IHDR   d   �   ��`
   	pHYs  D�  D�Z�H>   tEXtSoftware www.inkscape.org��<  |�IDATx��x�u6��lC$v��M�D��-[��ޔ��\�����s����%qI���%�ز�jJV/��E��c`��2�y�]��b�<���؝���sν�����|��?���4D�֛øL��0�����h#�G|�Ȉw�9�4��s"0�H4
˲��Iq;1���F`"�t�p�˄)��䙥���"���Ӧ��˲��{���Å7�E"��)�q��9�����0d2��`�p4\U����/Ek�O�[����0%��X/��֣�r�f�j�k���dĀð�2��0���Hx�i�-�y��K8>$�N�_S=�+��G��Z���+˲P����v?�wX����Jυ!X����7�y08�GR/I���{Q8�_f:V�6���/Ҝ�Q�:S�!�*�~���4��w��`�w.C��w+�#^���9�+�zPQ�����<���6қR蒭���� 0��V_�{g��i��yYB��>/��2�S��A��@h�u1>�aE53�C�6]c�˵pY.0<�lɱ0<\�o�o�@�$P� 2=P�jD��3��L��3��HH��S�(�� R=N��E:��JE���DPXXO�*d��`�PP�}|��?�����!��9[}ƀ�e�=�7�e��ro�	���4e}��d`�@�G���u�G��ZTfcԚ���S�i)N����F��I`HU�e��oDgG;��kp��!��c�
��ޏ��g�!F��2s&����������6:5c�/#�ӊ�"T�g (��0MDLַb\ĕ�L�s��L�p��q�'2�L7,O
֭�ɍ�`������I�?��St�Ěah����N��#��(u�Atx��!ܴu�N'�����L`�3���|I7�Ǧ>����b(�����v��������52��u+�������ԩiix����+@:Pe�V�c���1�r"g���R�C�{��=�����:ُ��V�Ǒ����ao|8繊X!S�\�_��Yz$���EX�0�=��K<"Ӄ������%�H�¬Lu�;��ڂ��f�fg�?P��A}���-��9s,1p23�`daR��is�K<:WC�~��� ��� ��+�B��ʩf�Q���Q?W�N,���(�0)�H�����g�8�,S"2K�x�:v��ظ���J�������R-~��o;_[�r-n}��Q��S�Ll�.�����EsaB�	5X��>���$1za�Į�6�������32���ya���<���Œd
m���ݸ��@���6�J�Y��q9PZ������2�SSSq�[�b�ǡ��YQ�{�2����ּ�����D9�֯���Fe�Y�N�!��5��N�sF���pj'nBTD�p,AF�ZDz�.� ׺*Q�D�M�t�{pߺ�9D��J�/�� ~��ӔW����&��om�B��'S���)�8����S)2+nӳE@(kʏR栬'��9��&43B���J�z9>���0eE�+F5C�l�.@S͸v�jB���n=�����Ӆ�HIq��%m��1��Fe�!�ȩ���x<���D�Ⴋ�n|��x��[9&�\�V<�f�芩�etQ���K��mK�wLM�ȼ��劝x>%�aaO3��ƭW](^� j[�f�,2�mX��?�zW���x�����RQ��ݽZd	c��b!���h'��q�=�k_�-�ZP{�#C�B8{�>7~�雒��~�ˤ�`n�7K�bn��cf���Dh�5Ob ���[���кu�mo��5�~F�`��o}��]�^�"�w�>'3�1�Ȓ��Զ�S��N�G�����aqQ����:"���h�i�����$�]#�k�E�
?
�{�o���7C���E��C�e���`�(��)���X����t}l�|7%?l�k+�,Ufո��@��}rN�M�}E��e��3�@�\g]&p|�)�Bw@��N��}~��/���P_��;?c(�2RR1un5:ח�_,}ŉ��"hP:{�a �B��w_�����������2j��Y
D=TXf���w!�`̡�����]|��6g��Br���V�Mlr�T}��zܑ�}��qи+��玅t�u��'�w �s��P��<�>��|�΅`)�h$xe�����yw�������p�2�,&��B�A�.G������r�@����v�KP��ϯ�a�Y�Q[�ޏ��L�t�Y)Z�#�m��ߺ���p�UR��VPB�c���}��)����BsW�2|J��nea�xŇIǑ��ro��o�Ȣ�r�h��3�����4�ۻA_嗡z�=*��ʈ�v	������ْ�Bbʈ�S���f˱��I
=���Os��ra��E<g��{B�%�y5��'�o�/г�Јf*g�:aD˘��=H8�F�g
cH-]}h��M:N]���Y�'״F��7#��'�*�Єt֕���LL�B6����N!;3C#BȈ��[~�t�lkC�&a��Z�#xܧő�����I�>�0R��q�[�2����aRӘ�G<?��E�-A5rW��&N2��n�H�F]�}�S��G	���ab����k42����~�GHTC��%�ʥDWbG���^Q����v8�M{i�>!���]'#��+d6쑁v����5Ƅ8�i��3�D�YL��+_ό��ےT=S��߯�)��'��ğ��%��ڜ��^-���J�}Q���ꁰoX�{a`A�5	�����/�CcS6oٍ~�睻�C^�'G�q��`^�h��Nq;7|�!�6y��ٚ��!��j=p��u�>Nf��k~n��n�C#�r5�ݟ:�N�X�rΔ��@o�nT�����E�3+ҵK�g$ch��5�[��|��}��f*}���
+���[n}:E���>��8�ԇg_> �ϯ�X��~�d�گ\�q������#zdS��!�k�H�D��i�VS�m)��H���|-�8;�Ӵ�ɿ)��d@�K��o)�3�أ��eT�C�Y�����\m����_`{�QQVQ�Sv��MF+�Jgs��?\ߊܜl���(&�R�I���3�������'��;��C#v�Be͵�`X�o�7h�Q3:^!sHx��wk��L�!@���z�Gϲ�1�H5)�Zk��[��ǖt��5ic�t�m��uԙ"qA��1���|˚v ��d�:�_Q���i�FCG�ٹii�����KǰqU)���o#8ѕ�={k�0����͸���$:��c��^�dN����}�`�$�P|8�D��@yn�C)��T���E)P�*�Xb�������Pb�/�8�A9�����Y�0Nߙz�L�sY�{Z�G����Tf�E2������F�Q�%�����Oh�o
����+3��˯Gfz:�{�/����y睏����;��/K�'PV����q��]���!�#�d�K�8�_���@�'��t���N"��RF�8��FL�ϴ��pb�@���G�!"Z�L���
WQ~�o�M��2�:���K�%�c���8g����C~CQ�,�}T�ɗ����Q��Lےm��6S9�-Q��~��aƙ5G����{0���k�Ava5z�|v�\�W^Qx�/�AE}�����!�[�FF�
���s�_�:�6+8�S.r9w���Q���� .k��SoAlؕ�utl�O�P�y�����(�E>=�k��`�c��p�8�qe�/���XzG��e��GQ-E��OZL�P�WD�4��&��.Mp��)�x��Y1o-J��+_�qآh��s��|�:kp��a!�$��A98SSR4M,mr�\���"����S���Q0�����7S2S��ze -�ax�p��S��'VGD�x�̊�#�R�T�c�����zݚ���>_�s��2��g��|㲨�ą�Z�cv�Z�����UQ�,�3���xQE��,����X�v�0�z�XZ�Z�碂|���`�;n/�F�_�߾�E��Iy��1\}���[���G:Dl���}�̎I�������!�P[�QX�Kh#��z��l�>,��x>�5.�q�UeЋ6qUqT���V������"��}˄�=�\��YE��i�oQ�SW�7�w|�QSb�e�ϳ��.n)��/�i���:2:C�V����\���bz�B0 �]Uj)ƿ2��٬�:�e��m���M�����2���Ey��"�a`ć���UV�̏��bi�M��WfQ���3�^����#p!8�C/��1�yy��j��v�DF��u!��j*P�h��C��ndF�ȧ��+#�:aB^O�X"�,�4q�0��g�𰥘��ce�:�D�M�!f���)KDZD���荠0���(�Ea?3`��e�GM�q?o�-��[�c(<�|�D�6 ��`
C2����Z	:�z����:����Z��1M<.Y����_Ӑ�8N��I^��R4Һ�����X�t$P��k?��9�Zy�R�����W��ֳ��c%$��C�u��}��>����˫�8C����]z�=ȷ g���}?^�DD�E�!���=��'�3���4�uΩ���p���a|y+Ѿ�
m�/��r�l��k;���i^�}�fh�}����i��st�����A�y�>��\=[|M}F#�w"�C�Q������u�ˬ�3(�X)"ks6D�w��3�Τ|��_\�w��Fj�<`�/����K��0$&f����	��]bu����"��1
��wdjǐ��2����溿�S��9��0^l~�2�Ǳ��{�rf���ç'Zw2M&�@��C��/N(	�t��/�I<��Q�0'�Wm��J�jI����*$abk�����~�ڦ�)�s���ul,L_Fkr��+��Q�,�9^��㽁9�N��8C ;gm5֯^	�o-M~lI=����g���zQ��Mg�w��yޟL��}4������d5KHG������{���Q��6���O��p����H������#�:�x&���3�������X]s����i��%�����B�A���<�0�(�������n�F�0��e]�ާ��e	v�a�h��8�֬ū����I�����dP�)�C��(�}t�~Ϊ��\����g�<�N�!�z��e�Ak$�/��@���c|�J~�N��1[�opE�`�m�z��~���{��{pϣ()Z���v\s�-C%#~�B��i��a<���u�����[���o':���p���8�=�v9��\&���j�>��C��5qa�^�]�pR��J��ݟ�݁L<�M�H<�e�����|�Y�����Kv�ɽ�P�6rr-��O�/@S��3�B����,��mmFv��DȇW�Q����8޲#]=�^������G1>95(�W�Sc�m�rY��CyӁ��q�w�"���y�D Y^V
����RGӢ�p��gb�7����)e['1dօ앸����z���C⪈4\�T��!����ӍVӊ�l���K0�ځg�]�2̆z׍��W����+�����I��|)$�ic^���)F�U�x��u���)�?�b���5ˀH����� �&3{浍���,�O�U8^����"��t��m?��I44w`�F Ý�����~����ՋUUh7#�GqC��𑵏#lD�]D�=�gɔ�p���J�>ӯ�j�hK��k�b�R�������@��*�~2�T���pݝ@��Y�w4���As<FqH0aH�i������w8/O#hn��YPR\�`I>*��HY�2W:��-�cA�����[�k���<�( �Y�8Ѯ�N��K�gT����$���a�py�!t{��4ߋ5�gEi�V���)�^���C�m���|�O��IhBz.(Љ=\%ܙ�A$�j���C���I��"Ί�v�i��LFo@	��?�}6�	�f��_�B���D�2���!p��HKq��H\�L�Bd�2�ϴ��qG̢����\òN�tN�il�%��B��䡉l�L�u�q��8��r$PW�x��Yz=�����dLGx�GGa#A3��OQ��c��+J���5Z��bw�q�E�Y�ь  �HF2�vT�C�5a��k�kx4 ��Y�ɥ_GO��HD-�(�g�Nn�F�TX{v��!"��'����X���24���c_A�Q�����b��س(�M@5�.тJ��`g��5�J)�&ų���d
gA<��"1��k�pџ5��>��v�߾^��`��I<����%�衮_S���A�#�]�'s�Ҕe��Z�ѷ(�ѹ9]����C�{��KPۥEӆ���e�un�1ad����D�aQ�)�$8�겁y҇k����E)b�8�vفh���[��_�~��6�
a��5�����f�e��ZQQ�oɰ��q͌�9Z����ז�O��FD���{S��l�bx���yE�e�:$C�l(Z�UL⡸$��:LAU-mP|�J'�<խgʩ����[/X4�lI~Hj��-p:~�I8*]mH+s��c^�Ta�(��xl0�Z[����S.,֩q��xM�r�����H�!ܔ�y���O���{R�\Z���uvj�v*3Ĵ�Фs��<U*��թ0 ��P��N�%CI��y8�IC��7mZ\P��3Wvc���g�	�i��GG:c\4h)Q�q��ӡ����,����6��'�:=.6�&m���N�����ֆÂ��1����&3n�p3
st�ӫ�mJ�l_]�|�a�$���a����X]F��Ɵ��ıƎS�MI��,����iZ�&<�^�"��e(���KD�M�25�����aŇ�t}NI����\r%��H�tK3-e9��I=#��#��P��Lv�=4��	�	O�M�k}��f�ZA\@�
�@hR�#y���<�h)Ԣw�w���(+)�������s�o��?�[�tܮ4d�`���H����4�!�`�ed�t#��!���o�V�����i�W�C��9�ۄJ�O2�\Uf0�k��o(e|Ǌ�B������TDq�k(3�2���&�%�rݖ��?hv(|/�d���M��c�jsVl����el�N���fBQ���{^��~���JI�����g�)�h�\z��AlX�k�_��6�����	7��f�4Xg�3�pN���Sk���LLa=҉!\>�=T,��p����Z?�VN�(��8��Æ��b@��>�������>��x�B$۔��.-O���,K� h��5�Q|@��!���f3�K���A��4�$5&�������I��-h'��w���>�b`h��l$N�N��r�jzz��#1MnٵQ��8�`k>�LӜ���BAT�����[r���oG��;�g�&&��D��Cs�����YQ
X-��VU�~gE��ho���d�YuSI�����X�OW$�o(�{����|��T��܋IC���2���v刓 [�`�ۻO��Q�e^VT�ʄ����E�X1���o(ǰ�Q�����.�S0j"�T���b�g�/ǊE�z��i�P�K<����h��܈�g����d�[��8�/�3i�����_�3��
Ky��E�l��P7f��C)ۿ]a)��P��y��E���`���`�Men��f��]��-�̽[�gM��/�uեbu�6j*k�#+-���R:�A;�;a�!�Q��s�������v��&�2��Z9�ҏ�T�b`�І�щ<E�@pJ�V /׸�Rp�bpkw�)�J���b5�u��O'BH_@�����}�0�[w�&��� [4"^}UiA��h*�0!���V�"A2���8��
�if�0!���Q��3P3(3Az��C�r�i�P!�i������"	�2�h}e�E�4��z�t��)aPD����D�s#AcVʳe:��{"LR��Jʹ����,���^-�,ģ�m����_�oB�VTZW�"N�!lӡc��]a��ψ2jd�#w��!,Wi���߀V��r�'+�����/|aB�(��嵓];/0l���`�AyU�����[m�u�ag��f�V��	k��I�^l�P�^]dQ����
��4i�����sŐP�`F%�R*lP2�ۛ5� ���9�pb�[5�4�� 4�
�R�*]�{�S;�$-q��Πf0@��=��3�,��=�>lz�'p�&��k)�9"�
���6��43�E�HB����(�z�	q�w1�N���:*@Pu�C;�]�$��� ��C�W��qLX�Jx����͈������b�Ո*;�fNq�o1id�W�&}�:�v�]��4.d����1C���rߨ�h\�`؝������i�J]�`k3j��3�P�Rlӥ5�	�()��s�`ṙ��(��2>]�8��{�"��g�W+9xZ�J�˥8t��aS��ljM��3�9��8N~��P�D�0�jI�NVUU��4$N`#��ո8�9�.ÊR?��	�o<k��P�C?'֡�p�'�ڎ<>�q��'�N�%AI�d%��q.v�a�(���M8^����Jdd��t�x��y?�95�0l3�?g�4�����W;=m�R�!g(o�Ɍ�G��1�Cc�'�=�g���[�Eė�x�Fd�#D������'^=��xekK��]�Do�ة��Q�����k�X����mL΃��sJ�F�f�0!�s�Rh�Sb��`�����xMuM�L�PK�d��-�hb���J�\�.���ʁ�[���:N�zV��;c��!�+�u%2�2��џY5�n�R{oT�"��#>��O����a�h�X���JEq:n�z;�<�����֚�u��5�abj/�<%(�)c{9#X'�7`)��Ԅz��Tx����xݒkS�������r���2+&�g|����w��:WZwn\����x����0CN�����A����G����%ȈX�����bez.�Bq(cT]����CDD�C�[t���qw��gXN��be�x��������j*��Xӄ0�����HM�V�
�s�� 7,a��Q	��$9��=ص�^	,��D��^^��ƾ��Sb�ti�������LW��3�����Ϣc$�@���L]��(��=2%8;x��K�EC!D&ŀ��(���][��{���ܵ�w�{��kzq*m�!&2�]�6I'Kp�}�Y���� r�}������D�L�Ҹ��X�Tb�hf��B�D"�-L���ܟ����f^��`D�<�
5��ĉ�L���TX��R���w�_����˥"s!��ŭ�~t?�Y9u?-�1�����`�9�hNk
��XS���M�"���v�
q�z����	�e�u�K�uĕ��e��d	���]bCw����A��i��@9�6,�ɿ��k���6/��,��*�k���aX���nꯗ1oc�.��-�PW��qw)����yHcE6w���IõW�2(���:���i5{���s1<�Ó�Ǉށ;R���^��߅uN]�B���:,N�:�8�Z�F�ԧ�s��2<���-22��$�k����Q�ߔ����;rm�{@�� ��x^�2d���p�E��z�L:s�%6�ך{���������{�cq��N�8`ffтD�R{AZ�ek�����F��ŹiB���ߏon���t-���%<��>�k�Nv�ͮ�K��M������Y��b�琨\{g��i��}�=�����9�d$C��A��y����N�+H�2z��E�5ˏ��0o3�"�;{�%�17�7=Sa��-Idq�O�s���
�V�M�0�P{�S�D#aXA��6��;�B��\�p�I9S�^`�^��ʑa^K���Zl���viq����q��D&���xQ�����6�AY�����hq�p����BYy���>8�.��<�@q�]ٚ��zs���h]��ݖ���Lʡ�!v�z�2�pO�~�QO�A�gNq���!;
�y�'#cDJrM�]��$�3�3�A=�8�_] ag���J��DK�}d~��@a-�92I�@"�@����\X��H3��:C�8*&Ἱ\+v��Ipvs�Fī"��z�	��e_y/�����d"H�2c�+u��!'Ӓw��ɬ�'��9�#�>1�SiI�^v &Kk���9m\-�<�'��Cv}yU(��߫�ր��(b8kHPދ��3I��֊��
�=|�}I��u*�%E���Q���S�0�2*}��s�j���Y����$bv M�����qD92��҅�C�I5�O�%c{5W��ִO1��
�&���"ai�RLQ�ƶ^��`�Gl���|Ƽ����X��G>˕%�<]��>{�
�����y���c��Zs���E�p��Mb�f��C0��"��ֵX^��fŉ�A����M+�q��m�z��o��e��R^8�c/���|�0�Yi�ӳ�6���s�xs�<��a��k?b8!<����#]��%rN������q�Nǘ~�,^��+�l�����>�M��a��1	�]��w��XGxr�]� &G�3@���,���H(��~�7���HOMŞ=���W_����*z<�aL�~Mu6��Y���_P&3���[�6=��z>������?ɘ�l�M���EX�����³�l����j���iʬ����(�ͱ�F�*���g4��>זFU�}V�n������urlW�� wv��w�Ԁj��y.KxĔ�:�>юT�?ou�k3���ԃ����ڡ�[߄Ԣ<tx���,[W�q�n3��Q|~?�;�Ԗw:M�>��@v�lm�2M�IX�������R�5�K��Fc��e��i��bexOUTm���^"��*��2��w�b���,<�c*�"E	�$�g	��^V	q��6�bX��mY����F/oZ,�YW�Kr���ˢj���5��(~�b�H4�зضq��C������U��g���*�3	��ii�j�Z'�{�.��`lA�t���f����rD�4����U>�6e�4f��@��e��Q���7��DuD�d��I����~�ͷ��'�ڼ�&)�A�;w�d	�+��h3�O��>Q����ʷR3�R#��"_��/�LU&�Y����37^YnÄ��WEGW�R��yy"����axF�93�������._��Q\w��x��oB �ï���*FQ��J�7�������0��^([V�PG���S>���*3j��q��Mݘ�U����u�s�"j�;�8?/��kP�Wei�?Yȑ�M�+����"{MT�h��}vm=�T��	�9/�R���,4�°K�0���CxqAT��8�w1�dY��f�P~��3%�.�N}�hl`$�34�+���J�{3�76�����d���8��08z�:���G��S�%���,�DX�B˶�g��A=nv́�ܐ����Gv��b�N��F�8����L�m�]v���*~�l��4��{�:���Cb���M|`�(��U�R	�O�vBx��P�2[Os�T�oo��}����b�ˁ;V�`��e��BV��p	Aы����d䩯���]�^?�FF�gV�c���t<���K���cW��V�l�+[�E-;f�?�RZL(G����w���G�-O�Wt<bu�~m��Ɑ��j�KqW�������9s:X��uGED�ڗYi[����!�o�0�Ym{�w�&w�򧄩���nOK��FZ�'_d&�u����__S�vB�oX�6ejLey&bJWY�;���$p_a�xźc�ym�L�H±Y�������5ȁ��]���o;s`kC{��=!�e���F�9]j<�"�9��%�M���?+H+���P�s�H��]7��Ș���5�����ܶT���%��\"~Hۄ(�,K�IVeX8���d<Cn�D�?��*��K��8�3���P�X�d~�X�Qo��&�+��ʯ8�Oc@�T��-�D��:�=iQB:������ĦU��_�U� �Rf�?��i�`K�l-s<j�#�Ĩ�x����=8���Hk"�+q6P4Y����V�L�a�glO�W�JQ4q֨��C���n��=w��;~�wm�x���������U#49�_�L`���Z�!/pT���g�S���c0(C/F���U�'����I�6���y�q�-́���I�����t�0)a��J���������܅s�߃�� jv�`!�q�bV��KOg��6�.Eu�G�O�
�����Jǁ�&�Gt�!ӱ� ���3�rPa�!���r�ڬt:���	8�ŋ^�O�aO&Ƈs�U�a,��;wo�u��S�]=��dDv�2���k��8w�6�t�܋/`���S�,ρxG^��8�Csf�R�e��c��K����ѱ�����9Y�������gams;�z�Ȝ��<�4셫ih��\�0�Ye��p���9�%C��9�<X?k�f3�23�[��_T��V���P�G��^��c<������:��4|��^��;�>a
�J2+Ob}���~��5+�W�ͷ�O��ڜ�Z�E�8�T��GqF�'(�����������T�!`��
���
N���-��/��XO難w8��u8�[:{�L�Ԗ��������v�����R޷���o��p8e����4��qE�c�:��˵��Q,�ƅ�I�aˊ�d�v.�u�����5�8�6���ϋ���-0�E�������|�?~�f���2�)��No�CXQ�(E��h kc�,�'��(�	M����9���s�=���^��$W���/��|^�TR�w}����Ť8S�,�ǲ�滆����ap*u�<Fc�q�03ص)�F�G�߃���q��x��ao@?�&��� F�	r�f=3QWߌ�^+�!��^j�pz�í�9�M��h������e͸�D��?g1<N�eg��������ڋ&���r4^|�2��=G�,�{�(ܬ
TP��9��EK-C���5���ح|s�r�,��-i��Q�OA^�r��-���Ox���HI�?w���UdUf��%Z\�~�aQ�e��LE�ŕ<"Eb`9���*�L�1�x{�6b�&���d�Lb�X�����e���9z2��aT�H��45���*؁y�DU�X��u�V��(9u�eW�X�@|�q�ɰ(���^�Ջpx"j��s�>Oe�2\wͥx��θ$?�أ��1��������Ȋ�P=�PBe됽T�rIY�NѢ"�A1;&�r-	G�┝QEൂ9����U��]�HT�m.����t����u-������ũ�l\&��׼�n*�-)�{�ޓ�����T�iSxgyZ�Ix�� 9J���\l޴{�������K�%��
LU����Xj�ոc��w,��Xi{��_S��n���͑M+�ˮ,K�m,�����L�E�
M�+쪤Sv	��	MX��>�������Mp6+^����-Xi�)�]f��b��
�KLM���T��9�z�j� ���kq�3_F�e�~�Ūp�[|��-p�1H�!r (3��W��,����:z�~#�j�*�������U+p"��U������l�e��n� �����X��לU-���:^Fa}��������f>I`���O<��D�)�Frde�+qC��%�d9Բ�B�OM�������'����ad����k�%�QU%4���W�����zy�Ojh�d��]yQ]�:������!S��ˊ�x~�TH��C��/��w��ˠ�<Kt����.p[
`�{_�UQ^b�؏t��/�5'�^���jJ<�9�ˊԖ�s��);�H���C�a��5�I���x�`5Ff�pTa#>����-D��PW}�V�$<�$��6����� ��FG�X�u�:�R;}��󺄤>4��d	%"��@�d�p�2K��0$b��d���).u3����厄��7�*��c�s��J�o���y�e����F�T
H����ˊ";+Mm�s.�'��)�h�x:�3��>å=�MK���̀�k�i$��|��۾a�/��0lj%���d.����@2��(�,��Fz�j{o�=��Y�)2;��k�|
3D%~f��ZIjOLN�D{���Fj�FԷvaR��9��U��܏����b R����L����$�>�����$��ek��q?Y?S�ߴ�!H1d�b^��lM"JX
��T��(����c�4�c����Z�r���f�[w����	�5�j���D C)����9}{AJ-Vq[�pf�,+F�kR#K�30��F�LˀD�W^\ ��n���`3���hh��'�t�p����ǯ���L/S���}����w�kJ�')�X���$1��hg�؞ٹ�O�S
"z1�����d�(K���a?�%�e��v�9u͔]�i׿�H�%�S�r�9��gѰUN+���\��J6����{cBF6��+�ބ��ו�������A�ç>#��(��׿�5��}.��oԹ#A`�Bi�r�e��2>��b�S<+�K���8�\�k�)>��5t����_i�z�����B�1�[�uf,}��m�ǘ��x��ޛ*�����eFo�Չ6w�$�_57WjB3�O��Q��L�a��O�5��v��"?٧�����EK��P�^a�}���ȼ�����,L
k���uk�zyjۇ��	Ŵ����1���J_'Q�J`���.�<)��de�:���}���5��,\]݁'~�p�NI�Ȥ�pT����
M z�Lڤ��!���z5<��߬�̬�Z!ؕ2�
���7Ӫ���I��c��W�5°ɵG�㨄&�Q�p���{d@���b��ш{��!�<O����SY-�5S9�Q)�Io��&����Ι�������Y��oۍx��g��%B�G��c�g1D�/Q.,�	�
�P�Dmc�
#��?>���h�߬4��Z�BSɫ~��,�f/�+���s���v��\�(7�i�#��4�|�Y(�e���w�)^�I�$����ig�X�X��b��H����(_^OF���5X���!�H_~�
t�/��Z�#u�:\{�[T���cM::������4S�vd֍U��۩��NdvU�.S�W�]=�k��dI��аkW���w�%x`�}(r}͡2��ی}�Im�z:q_���]�E�R$�"M z���Ә�8�=u�[�>+"�t���0���ø!Gg��Z�b���2Cn��C7�:�y���R��,T�H�-�\���$옌���G���[��չ����_��=Bȯ�������Ԭ��kR��7����ױ��\�+�f�*~�#��5�v(G�a���|#�*ߊ��ET~�'�6e���U�)sC#�L�����z���/���;�I��}z&�B�xY��E��|���H�����ɀ%���%wT�ssQ�o�Ժ�w�:�v]�>2��*x�
}uU̠����$�0-�gFs�����H���a���N$�f�3��FRVR�@%��Ire�x����3
�'D��`�2�"��ux�6�G]m3�{\����A�G�b�B9�k��{ �~��|N��������D�d	����u���f����s�D�'��O@��>.�Y���m���mL�;N|э�I�袠����5�2�%u�}ڣ�W����?���$w[�p�Y8܌{��3��Zꈽ7�9o�c��0X�<�������|�|�xID�ݳ33�J��w�m��ܕ����c(u�.<�:�l�yx�k�[u)궾f���\��b�QT��"�i�ߠA�TiU��Ж^�]d 1��i�3�9�%["���=���7UJ�Shb���q�p���Ȁs�U�X]�F�.�j���h��9]^I^Y�H��"�p#�����{��{�kߣ�.`C��'�=i6��d��u���]�k���C̌�6�T&���r�S�ħ�M�IB]�cTO�$�dl����T,|������e���x��T<]�ҫ�t
��T5.��b��f��I��*�`��#��!y#10�pmc���3ٸ�*�J�����{u��:���ׯ��u�0�׋��0�i�g|dÓpy�����xZ��n,�������ή =���CQ��K��b{JZx\��躳Q���7���i��P�a5�D�8]�D,��eE�w�8���Ĺ���t�s��*��xd7�F���P��5�/��ՙ��ܛ�]x�L<�b^�m����	�;%Ovv���b=֨|���<�ز����TU�f��K��A��"�<�h_���=���S�`�@��,�^c��3�-v�Mc�L�ێ��DǐX=\�N�����?K��b�|�ho�SJ�����B���`a�n�{k���_r���_��Q�����������?
���W]Y��j�p=ctԇ���xz��8���R�9�(5WS���^{�������&|���"r�s��>6�K�+]�p��bDCj	�@��;*�o�l�#���J9O�(&Z�bS�AQS[�5�����ƾg`ӎ��5_VUd#���ҒD��u��ԔT��*���*��5�{1�|~�f�AOp�аw��9[��YT��lMLCd�1�R�ކ�d�b��{�総��t�_��m�R��x�z��s��'���Rv��c׶�8��U��^RM�+��H)~IzZ*��d��7����t�vj�^�z~�U3�D+hY�o���]��0e� ��B���M��wV]�4�_r4�u�-z �jFx2�=a�ƙ��ݏ��LC���t�=w�z��@&�Aii)JT��9	=�E#�Y�]����ʝJO6�HE�7��(o��aN4�g��\�:������v��+��Dx���!�ŝ��?|_��ϕ�"�k���J�nV%6U�v�9�X\9��*�z����Y��0?
����G���YF��9������n�b���4���g�JX�}�*�p~��>t�'�,z�G�����ɨ傔oԏ�5'c����w����ձ��BY��Ѽ��H{1��,�̚�Мq�٥s�bc��8���oq�[S-�9#�EB�H���x�q,R&�#�?��o\`���j�E�V}C�WT(3����e��q�h�20f�W����1����ܘ~7�ҲpN�Z&~�P���;Y����'^�+\��ٜ����ם9 �)T���[w"%%��݇�Fې���x)rѬ�L͙���4w��x�_)��?b�p�����tt����a�蕃GeT�@���A_؅�U>Lչ�K�1��\mޮ�K�{�ڰ&��_�ԹLK�5g��\����h���B�Υ�B�uL�-��,�����yv!e�"�ކj����0��F�92 ��Z5���B��� ܸn�����ر�"t{'�Q�D��߲u���7K�j·~׵��X��Bq,�&�s��<ؽ�\44ԋ��G�F~���؉J�� vX{�ѱ$.Ѳ(�������^MX�2� ��̡��r+���Hh�9�F�b����в�)��n��b�:���	ꎕ/guR+x>�bᅘ�\��;��Ao��$7%��ߡ��/j�q���x��vn�G?�.|�?�C=��x�����9P��Ş~��C�(�V���?�^(g	���`�=��fi��{'�zM��'����R'��9�.�}pX�	gh��f��_M@����K�"2��W�1S�H�{B��f�/�G�0��52���c�5��,���,�y�����G�����р�y�萒������@e��y���@�ս�)�A�	4�ZĽmڬ�P�~..Y�	���eZ�n�Cs��-�h���`��a4��׎04A<E&S�1*�Xٖ�m�;?J��#�����z��a�Ⱂx7i=�Ul
G�6ގU��1"`�E����V�GNQ�|�bD>�@�~���"����yڛg�Ay��C��&�W��S�0����WP��e�q��9���,�̙Tk_�������l�Z�������ϭCb`kŌE*ԫ�����N��g�S��$J�0�N�1���_�������Tψ���oI8*�?��u�$�5��"���Q��5�5	�|�M�Ř:���~7u!f��&�\�w��yUV�*�S�sf���e;]s���֋w�]tŶ��i]�m���T�ؾS��Ch�Pϰ�8��dg	����s��f��6��$:t$6���(wj}T�pQZd�^�u��"]��s�+�``G۰E>���e��D{�ďذr�
�L����ޭ�����۹c>��;�_��b A��XX� �L\�b�a$��少|8�r0��'�c)����$7��9'lEKr`Qt&�{�k��fJ��6Ɗ�#���$����٢�eϧ�Z�9NV�̇~��%�y�u�G� �1Й���l7"�unyQ�:7�}y/&F��+�M���gc�;�P�\Ϛ��F|�����U����^��u$:�!����vIy�ܞ?����X���'T�ZZf��v��q�X��T%�'��O��P��b�D"Ac��$"��1�B��{Ėdy��,����!3R]z�	��V�~�Y �r�fD]�����<�<������wz)�BЯ~�߱r�r��}S���Z��"�$�y��{QD��x����R�I&�r�0�ͪl3U"�������2���JǗI����ߛ�E�djt���FtQ�����,�tUU�g����M�<w�!��-�mUZ�Qw��n���ʚz������*�BP�~����Y�e�\�+�xW��Ո��x�T9�sp/���a�5�;�7�͜dF���>���w���\��xD���ɩyv�o�R�&�qIƟE� ۘ��Qt�n�/T�z��E���]������:b��r�Sk�!�0&1���f-�iaQ�т�~��i�b���}a�
���*����Q�O�A�~���F�.����ǐ0��2��J��r�DV�)#�p�VDjV-��uW]��lqd$z�)x������a�����Ρ�;Q]U)��J��'��C#^��గǓJ�3�gUU�z�`�0b`��4��տ�BG:J\�GVh�4?z�XX�ztҹ��L��Tw�>-.z�i�x����g��<�R�2�Bk�{J1�a����������j�O�ի�g�
�k練(�]:��@o� *W�DZzں��'�Jas&���l��Z��u/���W^{�����!p ��u�fo��R���Y\���s�&���އ�~�'*���-�T�7�w��-ۤho]c���c���x&�s��4h�������zZ��h��'Vk"��cz#0�tΆ�ib��<��yZXT�\I�C�0��;w�~Y���LQD3�"�2[#�f@�D�0%��o��x`܋��E:�f9��y=u{��dչ(�����ߵ�����=O읎Z˛g��$]�����j�i+Z+�$��(�(��}��څa�7a'�D�䠽���TBpє�)����ƳC��ß2�=��k}���[b����ev<ܧ��!��A�#k�����?j���#�%��3$�m+��LF��T�� �p�q�2��?,����7U����ӽ}�v�8SXv���#��5�2�W���o۠�^'2��w��αB�s�ߑ0����5D�?�˘#�-�.-)��5딨:w�&�s�8�z�ժ�a��g��xK����aL��Ӊ��Z���3<`i{����-)��ϭ4�7'��1V�_.�١����!��I����?٫�M}�ml��[:���*��!kh���M����s��r:b3�C�5+[V'�p�d��R�)��#���W��u�Ƭ�7��A�0C%�8b���gM��Ȟ,�% ��is�8��}�M$�e��|�K0{��ji�^�'�J��cksv]L!O���>;I{���,����P^#<�u��Qw̵b8o�ͥ؅�	c�e�Z{�)5.�������ΟT�$t�]퇍~�w���+Ǉ�c���c3���|CXްF4r����"x`�|ù`E3���C.1�B�Ff�!��M굓�|�(���{ʹ�S�h0���AA��]��������t��k;�@
��l�0�R{P�{_�́���P)^,�&p���)5C[f��XƉf��m�.�䦒,<�<mz�O��8c���Ι�Hg��HG���Ś��<�5ܶ��մ����痟�Nq���no��L$|ɘ����ǚw�z�"̈�Nfz���r1�F3�n\�u���BC�2,�4�c�
/�:����,:�c:�`�̦��d�Cc�Z�gpf=���q*-aM=��o�=��z�a�؎绯�'�~��qǜ�c��;��VO{/�@��΍�QĪ�b��Ca0��W��u�K鰔��0�5b�`�N}�%,�B�/sW��'�}_�Y�	g1&ʮ�9��y;���l��?�K����(c�	����K�����_@a�Vۋ7��$ã8��91_�j�bf�SA�H�-��q#����Ϊu�N�c��\���� ���PG`ն�a{Kn�|U���Ofο����W��'0%�W��(^�k f�5��Ck�O>z?F|#�^�u{?z�V���ˇ����n�sa�7�:�������.�+�1�T��Mybe�$Kq������+�᪝��&���,�Hő���ft��,��ŔW@OZ��y$'�N����ᨵ���r��4-O�8X�Ͳ����.U�}<��I�v/�����~w*j䴔g}]Fr�C��t�4��o�Kl�8�:�
��t��n3�ZG��S_�kD��؀�����LN%��k��̸{9�����jv(�0��q�5�X��%�c���6�0jE\E0���@��ii�|��Ͳ�����$�	WՊ!ˍ�����,�}��8Z�%ĪJZ�t��6�NL �q=�@*�X��$��1�k�8�u���x��+�^"���h�>�x|��z7����+0�����_�g�R�T̿x� �SA�ff���S��M���g_=�)��Y�&U:r��+���NC�X?.�/\��7e���7���c����ubuc@��Cz��e�8���"��"�A@"C�V����~�$xl�n���C��b��y&���
���{��W�.���Ӑ���Zb��9��b�:��WQ��v��1��ۿ�֒�w]��s��'a���S�I�:K#>?\Nbw���h0��V��չ'�3�gj��K&��5���&cN\��&I Ƥ\ !�c�.$�'���ǖq)�L�b�&K��͠W	a%X����� ��8@�?�9\׌�ԔiO]�#"=��%qE��k�}Jc��N��_�W4�kuU%��;1�V������5O���yhʺ��Fu*s�$V��-v9�uv�}2� h�I�(ܖ��oc\5dIp���������僝�+��|�b�k<�/��N���2nɛQQ{��&� ��q�?�=G*	lM��ѺF��(@���g��FC��0�����`�רsI ��h�i�D����٬gь���6*�G����-GE����k4*c�y��I�3� o�S�3!�x;���D��l��{f�-n���ęmz��ʳ���==;d�gf�;����ۍJ����:�]a�D3����mH>+g����D�M S8C\�L�܏Enl=[3�BH��nj�lv�i�	��M�#u�@QsT�,z[�-�¶M�Te���.���y=u�f-q/n�D!ފ3���b�BZ]dEG0K,M�/�@�	C+	��RЖ�s�P!�F��bR��^
�(�_�L3���� ��"
�dEZ4^j�PP�D��ӆ�D�	眮���w�ȏ���y7=���t�ZD��/jFpA)�R�Њ"^����;%��Q�LaX�m��C������X������H|�M2�� ��ڑ�g�v")��b٥�Y����&&��7�ͫ�D��͆�.mI����8��Gp*-	���V�L�Ǳ��d�k��{�ɍ��biE���Gl�f�(f��L�;�}ּ��}]�ߑ��ÿ�������Y�dϰ�1}~]���5��i]�-#J�0ame	ʳL��D0>9�*�:R\���{�s�/.�m4!h�/z#�}/�^�䜣���BQ��?�@�r�!+��Ť��<-�|!�G8�'���߮�m�Jq��M=A��m�0B�B\{`�(� C���C$�M?�Ę��ִs�J"M-���a��8B2�R�RQP�V(��X�^2�;?�!N45���s
>Z[_���Ǹ���Q��ru�1�SmB4k����������I�z\��
��j�[������K*5��r!�G+N��1T�"�>�Z�t���o�W�J�`�h7pA�3���~X��R�L�1Աr�����i�ߏ�־
�X�� l�T�kG����t:;[��d�_̴��\x�N�����7�֬�B�Y�H�����1x�*5���[Ą��z>so�9��E�����<���Rl-�Ǫ�?"�^�o`�L<ۯ�ӗ SHTfQQ�����M&x�~k���L���oE��G$�C�$~{�&�7k���͙�{2�pR#��Q�@֌�����*!'�yy��?&bh��!��[~ݚ�(��Wq��FVf&���r�����I#d�%�='i�~�U�^Q�������֎�a@�p� J��ŉ1?�F
<��,�.c�\d�7�y�3!�ۄ ��Q+v��Te��_D�����b �o5hs�X`�'�ULgК���j�#��z�Y�˚�񤸢h�7OS�m'���Ch\��ۏ�e%p���76��"-ך���z?R�q�p�ZG.8#�mߩ
���W�4��w���P�\�v<�d|Z���YhhjEFzr�3����vJ���w��M��YAè�o?�h�7p�Z�����,p��<-Ǚ���E�7괉�<q��[���WCl�ֈw&��ƜZkL{��9�o[uz�yy:����eޥ��#'��V�Mk��8�.+ֺ��S��߿�\gg������t�Q}�j�3�54�GliikjG}{�=[�J�<��A}Q�X�Ǝt�F��1!����C�w	㯾��~��}p8�d���ڻ�8���]A�C/p�$vR$e��$J�DJ��HV,%q���Kv�e;ű'q���3qfܥȎU,;V�EU��$�fE� �{��p��Z����w�XL��3$���߻���{�_���IN,*o��p#���LE�H�mbP�3��>�����S<�����xf�ح?l%��:&>߫�,+N������M5$�?4��Ʒ��t\���:U�U,�Ʒ����ף]��UbC�������}��a�x���=D��MJ�5K�b>�a��^ٰ�]5j���NE bz��a߱-���G0)X#	���_j\6ٽ�!����Rp	��'H峤 {���y11�=�L�~*V����(lM!�ϯ^#@��?my�Vg��k~�V�j���gBs��&uo���M�l���R��mP��g	�?����J�e�G3�8��B�(��IvB �ݣ�BR��F�뾅K��/�:R��_[���S��l?��a��a�ոMH `.֧�����޷pǭ7ʪ�ĂY�ޱ+[Bx��1�R�`�EA���X'���u[�4�^�@�令�LQ挜7�k��al��o�x/O�w��>S�c���d���ᑘ�u�D��M�6ԧ_��<�s�M��qiH@坳�*�&�1��9�t�п%{躕=3�UF �g�_�.WU��h\�	0�N5�cʑ��8
��5A�:zDD�~�.���� ������|��J����P��,]"�
������e�~.jXt�P�P+��\?�r�t��F>$.�`gjcd_5�MRqZ�_$j]�i=�����]X�f8꾅/��~q��<�e(5.�ȰRyi�Ю���ED<m�;K�	���/59���xݕ ݤj-dƝ�nǚ���y�>�:�{���mBG~}���/Ǯ�}�)By�֍��O��� i��Fa�0���˅�N�-����h�I"�{L�2��1�hc�1���S��6�7_,����=��B�������]ې+4�����=�"X�_#.��X�p�2���g�&��]���h�z	�I����.櫮���y�nu���^{�/j��^zs�U���0G��2-���1<6)�U#jI��ГY�u�?lN�U����6����Mb���P�jǋs_���ׅ�V�֒������O��S����~ƺ&��"�f`j��7m���(j��P�W�A�x�IH-���b��n�\L9,]#b�Rr��s3��"�s��Ԟk��a��,��a��aαOͼ��S|,\P���[�EI����}s��wp���.���y(]Y*�LY�o~h�*������<�I��S\��=�$2rRq��7Bo௬p���8��i�_�B�aM�XDI\j<�t�-��e�?�y����%�F�_�����3�;�B6Yq '	>���P����Es��^�aIJ����n��D}?��PR�=�r�0��r�Ǌ��c{��c�Qb��!�l�M8,��@a�z�e�4|b+W�f��E��;O�ō��*�ʢ�>s��N���{�x敃Hΰ�C.J���Q/��-vnۂ���7��JC�Ƽ�ἅ��eLJ-MՅ�h�
bxP��t�
,�g~-��Un�O�7��e1~!V-�CW@j|�fJ��"3ۆ�!g�bp�{�AQA�l ɔ��-�*�%��n4t����)���)�s���"/���>[����ǓCm6:5�J�"�na7�Ǔ��T+n�v��ǰ��_ƟFh��o� 2�L�o? l�H�;�#eŅ�����V��#����!+�1��7����:>�:��
���AA��J�*\vhPU���Uj��w� FOi:N-]���Q���B�2*N>��S����X�R�>�{^�9v�=4�C��?���a��w�FhYda����2Y�IX�9�YX^�@M����l�ù�I�>o���fVh�?�ɺ��w��R�u9�(g�!3�	�_�%	�uKѻ��(mFu�jZ5��Ȳ��e�uB��,0O�#�3������0������Z����(�����\Y�.�sѤK��%��4�n�[]hh�De�$�;G���V�J�yy����9��auR@��T�N��Z�;Hjg�Jg�v+���<���5XɁȔ]���9��6�P4*�������|�T:�X���~�����6��SR������I���G���a�C[�x�l9�=������Tm}�"�*|v�EZ�w��B/�-/v~���]baN%ߍ��>�j\h
�j�B�sS\����C˓B/,��|�h�;�J0c�OuFƊ�t�wT#	'%�fT����$ k�wi�)]&��R�;+�%�kT��F�38� ��c�.���8�:^sN�]3*I�
Ń9A�`��_��&VW���c`����z!�r�-^����Z�zWio��!����k?�~t�T�P�x�R����N�A]͚S@���?�X�����V~�E�6�(~�F<�F�y���u�ߦxD	(�"?�k�>VE�C��[��#¹�o�vEȸZ��*ޡ/�ē�E�c�9����6�����/��/�v�.vL�e�����|�!fuz�����O���|�k�,#�ݪ��W�BA'�kP�(���/V����r�V.E��!�fe-��nfy�t(�a�9�K�k`���y=m�$R��Y��ɲ�!-	�&���D�Fx���aIb�
�P��[���5t�� ?�*�K�6F�] ��z�Y~x����2����]�݌�
��lc{r�F��	�BU��&p�,P�.C�DF��
��R�>�_%�0�tFW�&T�������6�M
�C�.ѥ�(����5����:'��(]��x�E���=�����s�$ɼKA�����N�l�>�ޘ,�����]���g��M��^,��!â/�1<�B�r������KْB��Yx$;w:ˁ�'�(��r���N�Ô4F�$k"��?I��gk�Zt�h97Һi�0P3#!7,�߲���&	�P/D��}ظb	6.+�aEG�0�Զ��k� ;+N���[�ܬ4�ؘ�υ��l��_7�Hb����!>��������&*`6�p�|�ZU�SeP��S�-rSX�����a-�j�:J��(���iե�M�*�BB��u�&�Ң�6��N�9y����4rU�7�Re�pO�IaE�س`MN	��)I��/���nڍ��t�9}o�}�V��-��(�>�l��!��ၹ���
�V+v�x���mEQA��=k��eES��f�>���#^�)a�W&n��B5��dA��
J�`�Ab�UY��(��̩�~'�(��F�/���@W/R�i�f[-Qv�O���;�~6?���} CO���������`Iu5څen��D����EO_?��~��զ�\x��)��磬`�4 �⃩t�">I��J�A���l��<o�,/�b�~K
RZ^�ߦ�=,�&<������4\�O�X}�p�i0��U>^��1��/t�gg	p���z��6���O��V�$ .�O�m��	F{�B��K���-2���� �-o�����L�Ҫ�ŰL��^q,��"S�v#��c@�������!g�W+@��\�ײsks��:��ֹ 6+��?}��>�,��<��;�O���G���H����5">�˙W��X�]+ң�
��-*�M6KV�Fe��д�)�?Z��D��}w�>Z�L=P+���� �����\���ԝU�������HG��+ĺſ>�y�줈�@�p/6_u�a��7
�##s�X�L�2�-�!ؘ9Xq��v�&U]�v�l����E.嵯^����hbYZ �*�hh��9#vJ�zF
YBs��ϫ�}���E"����v��\�`jb����YUJ���Z�)S�
t�KBХ?��)���FI�o�{?S��/Ԭ�B�I=T�-��΢� ��J����b��%B�շu�v��k�U$���O9161��6�ʿ�e���[�|c���'�# �G��K*�vu��M5$Nd�Ӛ�9�$�΅dG
ޘ�U=��K������ڂ�>��������?�*�}\��su&Ԟ^�^�o���pw3��,M�-Z�_Y!ܬ qTa���Wu~��L�#��jpݤ\S���Tɮ';��y%g�]�(l���)xyZ�#H9�l�r��ZG'��HM�=��x��~��+$7�֜���M�@$x;=�&��Y�BY� �e��'�BK���0]r3�;���@�4pN}y��0|�.Ӈ_������u*D�J�!]"\L��өX�!t��E{C����b��S��_�&����S*E�'oR�Ҥ�9����j>���4z�}�Of��<$TN��P{"����e��(�,z�)����m��U_��H�,�uL�'D�+�ZP�q�lGDL�/t�ZL=��8-�A�VuK�Kĵ�e6\mY��-����k�~u�FmP�ݢ���n����Oy+�lQ,o�H�o�xJ��9�^���Ţ���U����r�*��Y�ˁ�U����ꛇ���M�OHP�r��mYc���6��ͫ?$~������.�-�a��`w7BLi�����ӣ�*�	l�U�d�4���:�g���N�kǪ�?�la
�7c�5��ލ�Eym[Ƚg���s)p�\|�{@e��Vj�B���q��)d�'�0����VB��,��6a���	b�
��Y`Q�/ek��K+�ʾ��)��o�g�&T{cn��P�x��P��E#bw��%dG�b=T�����P���)��&��Pr�m?�sZ�2��]�־)p	�t���&��-;����/|�#x��}�rP��{b��S�"��~X��]̑�k�0I$S�8�Q���>ݹ�F"�@z��:���Q���1��x�EA��PSc��*�������
�醑��sk����T�O[����lb���n4\>1<���d,� ˜g,ħ�
�KuݢAmkp���1�G�+_e;'�C��p�5W���!��'�Ǳ�ވ��b!�\X=zL��7�rD}���`w�ar1;�G�\'k�+Q������HO��Ѻi`kW��|l�tR.��"ǡ ;3]��RS���ܞ� ���mx��Q�-�d=���ŧ��EF�-#Q�@�j0�eC��q��O/����e�0�׆k�n��� j�� /�C�M	��b5!���T_��}Ģ�,�����R���o��//���;�(��T�r�E{gO��!~��@?=�5K��ǆ�0>X���O�d�O�*�B?�A�s�}�['C��c�1�tb��ȫ*�ၬ�d|x�Z�9݉��$\���*s�ᣟ��fOuG�G+�^���f��'��2�*p���/m���L��`L142��I.O�Uu��qŎ9S 7�f���t�����d	-��� b��$(W����k�Z�uo���#�S��c��*s�������t9�ur�Gـ�y���"��i#��}��N��#\��~��A�P����I%蝝�As ��2�r��O��5�0�����W/�[r18����ā��K��dR.|��hY�y�T��1qt����M��rypŠ?b����N?�K�8�V9���?��ȼ!�oQNҳS14:3Oʪ�p~E���P�|���'ڃ��t�H{XZ�9$.��{~7kЪ���dŮ�kP���<����nDr�N7`�s~m�c��DM��q�q�d�-xQ4e���B�7hM+� @\b�>k���x�|�\`���U����ס{p #mH�,kbڃ��xD���`�C^=����y,뽎�j@&Y���d�P�����&�;h�����(B���b��"&���d��A�{�0E�AtRΰ�\�D14�(�K}!��-U���݃zN��n�U,ѡ�T���wͨ�H���Ĭ]W_��-9��U����"3*��V��5h�C�% ���I���kO�aT�׸{���A#@UQZ���\t��b��d���e�Q��x3T�T~�_Y�2r��pʥaUP�k	�\�W��tE�L��"��.�`G�����	.<��N�-8�S$ ���,%Ƅ��dS`B��9g��h�׵��(?���d|"�jG�@O�ټ[[��a����X�t��{�!�1��5E�׃%�NA}�SZ3�Q���3�v$��xl*�΀Q��9O�J����o.��$A�y:=�~(�6��ݳ¦�GL�9�ڠD��Ml58��"눎��㜄ţ	5���1��F�l��_>�dXĐ�{�/�Do��x)^���-�ehȿ�pT^+��#�Hc�C�R0��=��O�R�&1Fu}�jY6��zN���f}Ο��L�-�~�CH : 	Eb�x�˘	O��Z-].��{�B��Z�~E9R��8[�/�����:c�)�i�`�N�bL3 ��O.~��1�V��l����������\46|�.�}�ډ�@��&jk<!s:�Z&�I�������Ǘ�x�O��֤���z�/��/3���~�2�����y���ql����+�#9[	WBp(�����񒲄�~M�R�����J�^�3J�igO��R�S����WsR�𤰚�U��}����X��Z�H����5H����� AȮ6V/GCK�F�aΎB�G�I��D+f(v�܌��4��Q&p'S��I��AL.$��Ȝ��]���&�5�DQB�.�Cb|-�H-�B� �E��a,�b������,�LI
���,X��|GPN���.D�7B�I�A
M���2g!<,�_����X�w�#\t�e�P�r^jQ��D��d�>Y?�s��ei</�@$:���O��&�D P�w�f�2�[␆_k�0��k�m[V�rK4^=ր��ll_oĚA�H>����K��pKݸ�-ݱ@�7���ɷ����k;�V��� ��|�F��`̫����T��jy5�������b�a�8���!�Ip��f�E���c��O�'���BFz��s�¦��Fjnr2����fg�Q��M��x�λA45�,2��n���U*-�>,���+e���ʡH4�O˒�L�Q*�R�3�V�.&�)OS�:��D�0��0�K�o�a���t�A�.�6���|�MP�@�{����o148��;���t��G�jau��Ů��2���نTU-E^�Y�^��$��}�\�NH@�HK�BX�-u��;J�(c�vY�О��I�N�C����åJ]���ny�:K���-�_:��b�P2�%,?�ndi<a�r�h�vJ����^h����0%�>���+NǺ�*��W
�8���!���F���b��vئ�u�~=$ �aX	���yt��?Q2D�(�M�^�$,�,-�3�,u��ؕ��8F>���	�|��5�ւ�"�2�Dy�Y�&��dQ�}�G�?	e����-��}*˖��x��Aՙ�co�"P"�.%7���^/�'�:],�@ؚ��W��e	�vz�<؃�[�`����4��5]�ld�l@��s˽� PH���$	������n�^X��0K�Ȑׅj�*�§������.c��`���F� ��� 7�)�E.O��Z�W��,�&kvg�i/v�O����ʥ@ل)���P}� ��	��7l�R�K����~X���Ci�ӵ2�'�%��:5�&md��y6F�'P�����Mr���1���	�ְ�S�"k�{ܳd�c��]�Rov��1�/��~D^˅���<u:��xO�Jӫ3��FU�l��v����e�������
��Q�E���
0�ge������_�R�~� XW��tM�@���Ed:���b�e��\��[۲
B��-B��N�O�V����:�ѡ�I���Z.L�����.`�E��%Sh��;|{h�Eq,H�wʝ�kg���f�Z>J���\�H�|]��.�Vj�T	ا{��ĺ�$��5�E2�A,�w[�\��YU�4BFY����w*3&u���T�*1�,����#�{H�u�D�&A,@��+��I+�R�_�'����QhyE�1���8{�;�5�#���_�{s�s�!tH�{h��+�����3���]��C�D��*N���y2(��ߋ5�Ј��"Hq���P@�L�?1��,5x�墌��C~iK�%-�N��2��07�6�m6a�+,�w����*?�;Hx�iS}Ș���� Q���]���H�'c�X��4���q��RR��5%���(�����+��d����	��"(�TvG�]^�#���V�e��|L8�B�c��͞�[� �����I)v��ax��9/�\^���Ƌ���wplc�n􏊟c㘝���p���"d�8BYy��e���Y<��	��d!G�KUo�y�w����p:���ֈ²%�D�I��`Qq%�Xf��Pw��T�x0.�PY~/^���KzV���J����~YX���s�;6�g��ȃe<r9�bͅ��;e�?�W>|M>�f    IEND�B`�PK   ��X�z��kW S� /   images/65d233e5-7445-4b75-a6a5-2d8c2ad1af28.pngl\	8������)�6S�BDe�ci!{�K��c��j�1C��%{IY���14�>���,������:��L����r?�s?�7s]�Tݹ��v�v�]Rց����u�V��֭ߦ��6�ϫ�m�϶�X��9]��� �
��J=]��׋W]u�\1�]nAF���my�閘��uܘ�A:�)�������~�M6%1hSq�}��z�����H8{�YK�3�;gWF��~�J��L�<<b���FĶ�7����=�90�kD'��޺	�󗾝�|���o�{>��|*�H�3���F�)�> �l������v���9o�����ퟭ�՘ (a�S�@����(Y޼x_�fϚ���h��Y�C��5"0CB\5�[6FGn�`�z'�!���)����!���P&��{=9�Ȅ��p�c֟���|b���Q���2Z���&�쵭c��\.�Z&E�vx%ڳi�V��&�ua�d�x4�p���x���V�$�T2�8���`�I������O;`c��2큈�Hp��G:��m/�s�D��1��ڔ]�Y��&(ƌ2ܔ�"ʿ� _s����g��+�r����[}l����ۮ|{�`���}SsN��Y��^o��ꭖ��[�T�O܊
e�ڽl|��Cm	�	!��t;Vf �Lu�η��1Y?���R�>V��D�1AӬ�LPr��@M�77_!~3�;Ś�㦚��Sm���p䛐~�s�ř���Ե��4�uP��H�/2���˅���L��RC����	CT�ڭ�}�/V���H+ɍ	�Z����Y��q�o�X�%p��-�=Q~�1R�J �y�,	A�	w��o9`��~��,�k7�j?�2�����7��߼�x Y��&�1�j+�Dӟ���%�e{�%؍��_h���3�~�����h�f߂[e��ţ᠝с}|@�ȱ�!�������H���h���aMi8��'͜X��]5�<�ܔ�JUÆ�f�a��//<l�Gb>�P왺�}��W����M�X��9����^O��)�0N���E��a�X��jճ���t�,��q9����� }��"VW�8�ɖ��wn��"�}n�(O�F�	��掤P^��~�Ee�XTu�3��Z�z�s``���u��)Q�\�����"�ڝ�C/qS2=�F���SyZP���
G,YYȳɺ ]�c��lW�k�m�0�q(��B�!���u��R06��K����ГP�l�������w9x��1���1�6)買�ʧ�a�B��v�[83VB[�_�D
��d�z��	�;m`1fWB0ְ�Zޚ|��[�G:�`�L�4�� �/ԍOr�+�4a��l�$� �VvD�V.٩�(8��NX�q�r[F�W𣣣�1:�[a$Bh�vm��wZ^���dاo��˚̌хh���߷oI�l� ��_��*וv.�yqn��Z���7'$_���We��ٿԕ"����c���n�L���{Q�N�sPhg�����ъ���7*Gw��N#���]����w �^��_��|<�a�>!�#���Ѭ��-ܙ&���p��gL�n$�O��tN/c��C6�f �u �,h!�"��c�6ha����V]��-����WK���=1�-T���mE|��֌����v��Љ��Uv݈�؅�.�� �Y���0�r˺��l����@&oIcti1Y��b	!��.qGc-�_3�h5{%��k��3�ru�ϣ/���n'_�7t������7:N�ڭ�[ 	9��(!8V;����Q26�;) �J�7JF��%�6�@��{IFzVق�� z#H*#�*U���3@�1{����Lf��C�%��V�@����	s�}^�C�,`�gřZ�d~/{��S!a�6aq��L�A�=zF�
���r9&o`�� �ֱ���� k��{Y�v��(��9V�7 �"�Eא���u�?�d�m�!c���U���7�Q_����x�p���?����Q�[ܱ5���7,Q"<��+�p癁;O\��[����2A���U!���n����5�bת�B����s޺(2�oK,��T��b�����s^���� ��d���fH��U����8�ZÃY�����W����V\�����U�&�Z�_�����5�=hE.�����N;��TC����;�=�? ̲cs9r�6
-;�J�3dHN�;S���_�������3h8���e
v��%B�HtCV9ޛW�k��ǰY#�%�
�w�6����Yiw�<O\����t����M�ν�7��+P���h����[�1D&��t&�{�A��f�4�+�16�O���tQZ�K+O�ii7[�#�d�3��Oe�f�oT� ��.V	�%��Uh'����=Wq�f�Ww�."
[8&.ʒ9����[�KtQ;8��-O���h�ٞ������-�X�z=�{�d�z,N�$��6�@q��r��R�ws�?�Y��0_)B`­$�8����}�o�no!��1�j���3GG�����s����(���9�/�6ǜA��9��5� g	ģ<�\v�By�:��,Kf���/OKcg��$�9yӴ�cNě���;�7"K��Ey��	���h��H胈Z����n]�����G5|��#�m�-�uQ���O�ޗP�p�UY߅釨�
�=�t�#޽�^��*B�j�-�7��!�R���R��to�\��8�;La6&y��@@�@��*!�U��p�S9��%N ����	-�8/�i�Ä���9�������Y^��	�V�.4g��E�\�0m.��X�W���w�=2����>�_���N ��(
A��RUϑ���	56vw�|��%�a�B,-?Q�'-��DD3�*�G��!�{M�g��g��Y� ��k���x����!N��#�*�1SZ_�ZM__[_��
�5>��M���`1y]T����O�Bz��?d]Kz����"=A/�rL�q8�?��uBǞ�G��,�*�̴�;v�{��bf�U+� c]�N�+p$-Ge���h񹀢d� �h
��]���&�B�(J-n�ĥ���"+.O����a�g��}��Ytt�!�h�s���3�\[!x3&�����&�<[�\�T����{���)N<�����uK��"E��̵�<��$�y��I�w �yԀ���f�z">�yJ'&R;�ptmf����*�:��c#�d�H�8mb�~~ϵV�*������=�666�(~6Pa7�������p(�����h�.�zJ�u����6��D�#�����/��S��8u:$���S�W��wq8ʢ��d=�{���5?����@�3�3����"D�Z׆��<��N(�^üu#��7��u�0�愸�9I��G��Y�+;�G~
7�"5�#{]G����y��+�xBuHJ�A/���J����!�	���"���������޻�7��.�͗�]��9Z�#��a��a�����O2.V�_���� �V�%�H���ח�ii#]�H�N��@����6_	~����y��_TQJ�������9������l�`�3:;����(5�mϟ
keF��
~x`G]]]�jUnjT���J����0�*-}}��T��rWVD��G{�����
,.YZ"���s���y�����S���C�cMX~�ݐ���+�᦯O���)peO!s�,�+��^��$��߶��	�;Ԧ��'|f�Br&����s}5�5��{���-,�����wT�
mVxz��͑p��N�f�8Mc�����"�70(��F��sJ"O,�$ڛ��2!hEl����z0�F���.e� o"��ҧ%%�i�r�3�W"/�a�{Ԣ)�ę����~A&r 쫗ݤ8�������˺2�-Mx�.;��������#&�j�Oo](�M���ɽ&����Sf�s�?䈷�;����W0���=�zy8��
hH���=����
�"�P����x���3ř!Lۥ�Mg�n�5�a���XG�@|rbFA=Trf��Q�+�D"<"n�����5��+�srHh��490H�*-0�HYn�}w4֕�ڧ�������f���Q!'�Y	��9B^��0[<�����m�]�%��%/��U�WxY�bǉ̜��lO��~1��;��h)/�`;L��M�s��hfV,���`���e�����Ak�o�	7Ŏ���c&�
���/&#M� ���"ZvE��L��!��?e��n�t\�<q�8�ۜ�ci�e��vFx��|��1�ʡ�}S.@0�(�<`��b��6+$�;�s�6��Pk��jQ:���e��61��dW���4S�t��f�`%fL|ˏʇ�f�3�ɑ�='E5Z�M۷R!����e`�UՒ��H!�N������uۀ����N��x�� ��U��@y�]xƊ�uk����~�1((��;�5�[#�YF���Ў�|�����������;���и���R����sӌ�׶$'&b�p�8�zJ�҆]���JKkV���3��N��/�4��~t@=X�3�c�xyP�+�bk�X�ױ(w(>��x��_,��q����ZU�;T�D'��,�[ǔ��:��R.<�6F��C�3`��L���C�����z|7�I��s�ʷ_����Q�B_g���u�"vI�ǆ����ol�(�?܋�'쥺{�T���|y.�(�s^v��g�:��A�,����b��h�Dw(��?���C��L�y1� }�@/��S|?ĺO����i��'����C(�IZ�M�W*��Ͳ��mP�+g�^S8-M��m�"�/�G͒v��!�u��*��Q�����$��i;t1g�y	��g����0�0x�E�y�\�"���(�}��6�J��vnE��: 雰�y�u�ף�בPpğm2*R��5���&i2Sc�+�Q%����y�Em`��r�YS��qX���Է�
d9� �?����(++�W-eT����x�� XZZ��EFr�:��BLb/<d[jMKŖ���*,�8���)"��WF��c�a)�8;$S>oB������A��:K�P⭟�C+,v����Hr��%�B:nP���Yx̠k���+S��Oz,?{��l?F��0���FKUg��77Y2��? �ܪ����;�T���Tai݀���� �������zIϲ0�>���g��\��,��_Tg�L<c�g$	H{�ª=@��Z7���we5�&�>561񹈢db���O4
��������K�؈T>4�:--��M��N����VP�^Ɣ]b��e׉_ ��ř�d���a����a~�`�?�~�8a/�"HX��p<�a�%��Be�� X�Z��~�562Z���b�>4�HȰ�M1�c	�����m��^��p��U�'����3%�\c�"B�m{�$��vԘgqq&��r�8~���UNs>�?e0Ն�rs`����?ղdwo�����N�\�T^�j>�e�������~��=�����/��uD�ꯂ�n#�����zOds �� �X,mTD����Dl��2Lj�Dj��T��iY�x���l���E���~��E_��̑T�dt횧#�7��c��x0�����Sü�Y���N%��b�ʣ⷏f�du\��1x<O�Koe��$��_����6?�����eW.Ã�3,��dd\\��?�MH%�Iu����>-敔��t�6�|�'Ӏ)���,vqL$��w6Kʒ�錦љW�� ���)��g)D]`r��"~��[���^⤡�|�'α���|%/˗��GbĢ��=+|�aܿZBO�}��zU��_����eR;�7�c��J|�����/_.�C�f�p`<$\�?����2bθm�ߕ�e��YH`��m�bq�O}lsE_�5�E��cBX�0ؒ��b@���
\%))8���ZJ ��ڃffܲ�%��F�\[' ��[=	]~�C�n|=*���8-5d�-�ie�|�'~�gwP��3�N$flњc�A�*A�j�n��{�O����Ihhx�[�!�������̒�� #yfa�z��K���t5�0��UNY��(T}�1Xm3�RR{D��eWg���T.c�o�n�t
:P� Q��5`:�O�>�A��yj �sDjY���ga�B= B�\?99Y@Ƒ�9JԻI��^�W���p�G�!�?��q��F�G��T+ ��4QЮ³O�`h�J�׮�gٔ��-s���~��@^ǣ��  �=B&K@����m.�e��^��Vr��d���e�̒�οbNn㲰�����Q"�𥳐�LkFF�8������r��Hl�����p<��M:L-��U��������\i�B^�f��J����7����ŵ�������7m'����N�*�1�;��nO�@�&}E��Zt�?K�u��ϧZ�^�F�ߴ�Y�z�e�x�Y���K�4�#'�޶�)�3L}��.v���,i]9f��ȴ]��MO?�)��Q����U@+�z�F�]8��f:�U33������C��Vp�'Nf�����" ��+�4 ��Ox�mX pÓT��gr�R�j�(d74���`;����䕒h�ߢ 	�?�9��9
<K��<E�y�Tb��l/��.B����Ɉ��4�^"X���#�i����Ȱ��"�Յף&O �j,$�♠8�0�����P*�e̶�x�JKC޻�(d?F�4Ѝ�<��fmڞ��f�jeΟV&���$$�>����q� �����@y�ׂEw(4��^������<����I���4��th�[�ŧnU�r����v�rl�Cv�}�Q9/���c��5�vq�AYrH�lzZ�W{E �c������-�z��X������*���b��Ye�G�D]��}~
��t��c��4Sr��:���h@����ZE\:y\L�OE��q�fw�����Y�R����bzT�vr�/<�<:�/�7��
� @�:=R�i�	�D'0�b�+�
�S*!],`d�*}=��͐��w'�ș�׮�>h�b�E >9 4R�(�N=0Z��}���z��y=�+���zZ;��6S�����C2gff�g��Ѽ3��D�*��U%�ޒ�=�A������	�_�a�"O�_�R�C��r�!��O�$��� 
����,,D6�prt�xj5���ȣm��:��z$����ֹ�O���Q��L����G�bۻ� q��Ro�[���߆Wf

*�ӟ�P6Q��=R�ڪ_��D�R���2�G�6��Fu� ����;�DibMC��(��3.+�ҩ]t�cǎ�+}�{��}>�9�lw`P��3�d�϶�ň�[�~���{�h��a<'��u�]����Y+�T���0��Gq�	���xeX����ҵ�'N��\���T�Td���n����BP�i$����Y�ӵ�q����y8�g � U��"�ٶ���?{�%��A���鍖666��~b�3Q� ��Mf&HWb�&h�fʞv3o��rԶu�$�亮Bd���%=����q�1f�����}�EJ��t���¹Ǒ͗j�`CC�|�1(@+=Mt�bm���_)!> e`�v�m��7~����u��ŪIC�A��Jv�E%�Z�[�3�`�o����!���
0�}4d�����=(a�٢S��SFI��S��^�Dt&�f�&BHyo�N�$ߔ:��;88X��Q���0d��(�D9^h���;������x~~�c�VX � !��pt�A�>��ISjZZ	h��C���u��:,��$�a���D:�I�SE�&&���2_o�����q	̫W��4�'0���ȧ�SGȠ�xa�n��ׁB�*��.� .�Ru�e���4������G�uhoT�E���c"$q�+{Ko���(�4w떸�K��I��x���	L/�>PQ};���Cl�J���w����pW\h
�~��x�/Ի��@���,�U�顴�(IG�8�(կ������g�^���
zh!t�Jz�����`Hw0�6�����A�%& \,���8�H��h��L^���iL�]�.<�Vv����ż�<�>�gBs�@O�د'd	l� �3Y0�����u�J؈���L�-=����E��.j����Z��ǣ��&]�Y?���̍���������"e��n@P*�A��a+�@��g��g��
�Wxg8��;��9~66F7g`{G������y|F���b�@��ü�}�hT]�<�%�q�܊C�c[���!��x=�۹�W�>;l+_�o�u�Aj�����{`�9�T��z�XO	}�[��k���쎎�6�á��qa�b+6�bz ����l�.�}����E���x��e�?G��?^��W?X����>ZE�bOT�d�^55�MI�m�����v�&��5��j�b;�������0��0z��i�O���
�����>g�}���,l���!&}%�泇3���z�7z�����>Pw��o!�T�l���*?��cϴP��� ���*�J8���D>֣I�����x
B����N۬�]���X��[=Wq���>�[�h_�2�+�z�H��>p����@;�?�/|>,���;��4���H�|;����X�VVɿ�;9�I(z8٢���M4v߇˜�=-���s��}e�k�a����-�2�Ehkߙ��y>UTTs��	J ��������MoRb�b��܏�$�/jj��V�ɡ$�E
N���<��K^;�����T	{�"�P�M_�GEE���^�G�!���1KMd)�����
]i��6�IW'�����Yp�d�����'hA�h4������8y�L�|=�,�B�G®�c���b���ހ;t�u��Ç{/C��F\�r��c05�1�&+�}�SQds* �q֩����t���oEig.�F�}�P��j�:-�8�]�j} ��S__�q�y�k��\�����3�]Kz4���cZ�������E���� �D���+�59��_�9�,�_�`g`�A�^�4�q��>DL�]F��\8�R���	O�o&f���m���I�f@��2�����a�����0740�=�v���[�f���	!�����s|4H�{���y��:�q���)N�d?P�|�)77L�RoA+��π���\E����z�F3rE+2� =���xv�8�k�{gA���/jK�ƭ5M�ڥ�>��?])����� �Rp�p�:��$���q
�G?�xX�覶������]�����<��#�{ە��w����U�}Pw�cţ��N/Y��F<X�v�������:*g�і���G40�zz Fe۔���4b��\5{L�VQ��4(�N__��� 	$��u��C�/'�n��ID&_Fە^�*��"3����;�y�����CJU���n����P5�_x={N� ���.$7��9n�Z!j�����܄���Hf:���b�]d�Հ��e�G����μc�̵Q��K��`���Y�K�������0���'��n�	]��M�M��ˑ̐�sX��Am�4.K!%F��18"���<�,�عj)�E���13�`̆b�؝��b%X$%@HJܩ�9%Z{KݎTV
X�2!�ݓ�\��B��c�[�[�Ѹ;}���X�f� L��Iu[�5�y��NM(O��h\�Q@��uLQ���
P�?�欄��/#:�K�X�}�Bq�r*�&�N��Fχ�?vw�X.2�x�lx0���_{���ԝ���o`1�O�+fʿ�#�k����!��%��y�f\�r���y��\%_�ڐ�k! �c
C�n���������i(y>Y�?�� P@IIl�,:8��i�FR�C͇�މ��n	x�fa0o�®��3��L��fD`����!�J"���b�%�F�;I������[��r/�9�<����Cӊ_���I�^�Lm�h�7��qn֭�,>�[�E�'Y�V�P�>�?����e	��Vd�����q�	���B4N�wA�A�);���o@-����B7��h�E6P/@��;�s��q���*�/y@x���t�rb�Ū�̟�@Á���E~P��x��M���s+�K�$j'��	$Y��Oo>w�f��?�q�omm��9Ùw^x�y��f;�s<W,x}�j#(�������P{��������K9q�y~o�:kIS׎2~C^���e^~������8�}��%����sU����Y��XW���nzy���/iG!(� ����?_�T������CqV---��3˯��ݼ�U_Z�~�ԃ���x4)e��$��t{8\�7݀���z��F|�U��t�c��O�ə�g5���J;�)�Z~�(�{�*���B��e�F�a�rZoKﭙ�ds֗�/ϘRw���~�>��6s�5�5J\�u�d	2TL���}}��5Ȟ:����VW�8���ɼ�1-?�.�g~P�޶�K�.�
_//92�q���!�,+��NP|��iW�/�2���pnj�Ƞ�,I^�A��N�5%DrʧO���?���7w��SW�����GԚ+����h���Y���^{��e��pb-��Nc\�)V'�̊j��*���;���NAX*��t�/�[=%8 �;��MK�쬍��g������M��N�y�8uܵ;��'�J�;�-~��0�_�e�}��<o<�UDa����70:��>"EБs�X�,C%�}A	�M�v+�͗�I�(���Y�Y��T��A>�=`�:��0�����+>IG䀥^V��*dq����YF᎕E���BJ�4A|�B��3�]6M��`-�<�j��x��=t!0̽�Q�!����$?�a�f��T�Nj���v%$��M-�VVw���D�Su��W�g�/�@Pcrr���
��"����}ư�6�1Z��&i��S�̄�='���~�5v5��HkMá}/+:�����_�q��bRۭ0���m!tD�*�w��{�V/3�êJ^�YRy�&g�"~�nj<�]GRҵX b��Ǒ�V`|�G~u�?��s���2�{^��y����5��i���U�ʳ+�m�@��f�Q'NW,U=�ӎ*N�c��2�0H����zuTG,z���!�"BP;�hf�Ң4S�joo�%�͵;.u�Y�y��LPivLr`���W�G���37&7]�ڵufl���Sa���$�_�Jd�Ȍ���>D�ĒK�[�h��V���v�Μ�-���17r7��;�ſ�?πa���E�,=��^�N��1.1s���S�g֬+�@�����S�:�5w�z~-|���_�+m�ś�(����<��%�-��d��S1Nlz��X¡˽*w��]�e�[b��� ���|���-K /�>c����8/��1����^^�5���M�~�t)��X_�D�����i�ׂjz��g�7s�tR51��Wñ�3;N���Ü�'w� I,���˫UW-o陭r^�-�[���X꟞�B���5�3ҏ�E��~ﯱȐ���*�ݢ�^k�u(|���E�VX����8c��iz�~y&�B�'�(�/}�L�)!>�L4t ��炒�<0��^�7|��mx+X��'�����cE�
Ki{��5K����r�l�����ռ����d,�Mk�����F��R���=&�5��̝n�>#���_B��B|����j.���"��Nȫ�ݚ��Ԭ=ݕ>�rGAlA1��Cj!*�4�k�2df��}��ǘ�>RZ��7��*����	�j��1�����T�-t1�V5ﮞ��r��>r�[��&��m
@����=�"0d� ��jg�����¡��Gy����S�2$U5�lo�����Tҝ�HA5�W�}�"�������t1��qݥO�S��ӮG)�TN7��/7��10�`����l����իJ�gz*��<)�]�o��ȼ�v�����m[p�m�w67�W-=��o�����?��ѴC��ƿL�B�s(���8`^��M����%���A�/��@4Ro=��ߝ�g�����M����^!��;y73콽m�\��
��8+]k�/�}X���ۉb��G�m��e@*gF��x��E$DEޱ�:%����Ö��?�
�,K`��a���:��Lj��{���MW��p��fs�&�Q�m<��3-.��/-h�z��K�ݭ���s�RK�+�����С���.>}��Z�	
W��$��c��P)-�����'��>˒��[G2��AlCm�;���g����2���U�a��B� �*y��M�{�.~��I�i$03��;�?�����Mp�����p%�L�ys��V�#K�a����� ��(5��~	�.��0�-���P��RO�����A�S�,ph%R�{��G8�6��r�A�~��h��vm`sb  U� �q^4j�g=���vϮ߀E!���Lu�Sգ��iY��SA�����ˎ@� 9.�o�d$�	t]~����]@�m����ʯ�n�5^wP-��2E}����S���c]��W ������0p�"�ĉ��ލ���/uL� �,��C�]+�'oԼ�Ez�:�ʢQ�wJ����]W�,ǡ�ns*X���Z��]�vIX k\�NMh�z7�%J5�|��Ӑ%�O�M,.���� ٟ�߃p�����,4����p~�F*^>��^C�P��ϔi5?��G�����@v�ךK#�NU㞺j6˒�-�cj�h���*�ߞZ^��3^*(�1�2Y�ZY0޵��Gk=�扈?.�ݺ"1�x�?�RT���sUO?6����@v���;�~��ʚ���/��֭�!*��5�r{:ְH��Vc��P,9�dK5"��X?
<��?I������ޡO���?�b��N�CC�RDf��e�����@�������\��Rw"�}J��YK��	��\��*f��KŪ���e{7W��[M�NMM��Th+�4-d_��!��>}�ܝ+�`�\��	t��.�(c����X$
_�{��i�ڮD>� �P� W��e�<.��eٝ�R����wD7�3�7�;�'(Bf~��}�gl�u�iA
�\��v@jyF��b��#��y��=�Z�3�j�w�@M�2ҒJ�%�L��?p���=�v%�h�x4����܌<%AJ����}N�O�俻]�2n��	@T<3A�_vb٪�ksg	&k����?p-���")�9��؂��"w�P�R��i	�M>���܇�f�Y:�i�s��A�S��V�u5Ev��^'�ǘ�(�]�5UP�A�x�4JV�x�P�l��}w�[�Ơ�����G-)ZJ?�_5�e]w5jF������0;�ڇ��1�+�z�a������W���D�=������۷��^'��㡖��je�[t�XT�'�ɒQ@�ڝV�RRR�Vw���+�m�u�<�Z�LU$2�t�$����͍����k��Z�V��u9p���-Ч���Js=�����PV�yaV<woP��qepnb�9r�y��
�hq��/��;�g��D�S[��>b~Q��uzX�eG��w�c����ǀ�Ů����GHZ�y���w��/�J��h����c��Zӆ"N.�P$9�ҍ���֩z�y��uF����^�D�M�s0���7����z;�[��E�H���;y�'0=n���e�N�;I��s�XkD	��Pf�6����zc�_�>Lq�5x�]���l��)�5�%���Ji�A6_�^T��X~e"�_�A�ð讪�Ҷ��Kzq5�Ѹz��}�wCG /��Roݐ+,_��]��H%QQ���"�%z�7�82�`�N����J��YNKII�t<�Y�������O��e�*�:�俲��)d<�m����!]x��� -S�s���9!Xr%Lr(�F'�y��r+���������Hϡ�{����^:�Wc�4��!\3�r��K�}�Fz��Pg��$����ч��ʆ�_�̝�J��˹��3a�[�C�;�-HEU1!���49y���{x�E��u*&��BP-R��(��O�J��KccM�δ�߿_T��he��?�>'jK�9�:^i�~&�@A�v�/!)t�����ۈ���F�!&5C�<��.�d\�l�,�K)%U��(�#��3MOtƈ�]5��Cf��1���g�¥�B�]a��˘>6�g���BSw ��W���>���5��a5{�x�f����D�//9��W��:e.�%�y�wTf���+�������_7ȳtAι�*�R,�NܙP��V9���b#��7;��q�M
�����)f�Q�ˈ�E��ϼ:�"���5��Q�rb�'>�K�4V���hm�X1�x���hy�m��AK? ���w�=�m���&k5����K��B���(�Se�Y~���S ���E���bQ�V.���*�"��Q˝����E�H�����O�O������u���]	�{,���._���I������f��E�Sd���6_���!��?!���)�q�%�o���e2)�J��-r�K��B~�����Gi�C�y��z�<V��
^��I�K^/iǉ�]�p	�.�xh�n;$������K����|��_G_�1��^�"�'-�v��3EQ0�v�!�|ya�:� 啘��&Vi����b:�@�_���[=y�G[t&�e��N�}ɢ�]-X[B&��f�u��K3⧫�_hF�Z3U�jn���ǯ49#���G�W�|�+4�R �B}�잵ʬk&����B������Hr��k=Q���1��W��Ay��E�����/ ��rg

�c,�3mZy���5�f�;�[LK�L�.�H�M��U.���B~�d?`i&BQ$yBﲮ_M����@&٣:@V�]��7r>m�!�6"�>�-^��b�����F+����T��d��N}3{#��۠23�,9�������S�xB�s��.��0��5�e�}�3�D}-n�,	�t|��'rW@Ơ�,|p��7�@B��Y��}�w���u�����$m�.S���̭T
�9��~���=O'U�gs��B�ZV�Q���A�k#�A5��;q��3U�ġǬ�nv�1�3�
���Q�{j&Z��~�����σ.�4��j�QT���-�6`�
����N�Oa���������}'�T6>��S#����!"c���\Y���: k���8�I�i	��Cɡ����W|�jز�Z� ��F��ދ��m����?�N1C�?�Uy�K�H.q�~JL�	0vN����k��.?�rQ�݀Z�7Uw^��*�����4ӮT���0�"w|�1��W��4�Q�<�^cc{�$ɿ�5�c��R��!��q�I�¶{)�^a�*>�ⷜ;[�e[�2KB�D�86��bY�,QI����r�9�<A�3�D�\�Y]���d���r�"i��ܞ����P���ѽ���~t���000����8`�l����s<�t���X_~�9� ��,��Sշ]\\��'!�v�m	$?7E@��,�O��'..6ׯ�ksP�<�k쬹Ob�)y��9G�	�~�[Η�"]�wX!�`.�q�z&�+�gvto蝧.%U���wz�K���Mz�z˝�)n5�1��P��Aw謖��S�1��.(`!!���\�|O��>Sm���stR#%��E�',oa}m_<X��jh�=�$1�a5��{���C�����5U7x��~wC�Cx�c�$6���~���l����>���[H��9G)3 �Q�.�Ĵa�^,���#� sz�]��9k�"�KVa�4�'��J�ti��GE���<��a�X�\�
�H��ĈK��w� &�@P���ͬ{�\��l;�-��.~��QhA�R_߃��1"Y.��؃�yjvy�M`����---Z�-��2,�!�˪)i�Ek1�6���lN�Ѥ���K��Td2���By��㫇ʀ5�V���!L�Uy��2899��IcvdLBN�e���( |�,�2̵�í�#��RԻF����zw҃�p�C�|�Ty;�O�8�T&���� �H�1���<�pjBԴ��aYɦ����`���J�K�و�G���[�w�E��RA[� ���ـ��:F1����s���{��s��Ӣ��w���sSw����0��cv����l(����oAl9���������s��h���,�?(�E$���B�7�m�R��W���!����C�T��vөCۊ�
�쵝���>��E�)9�U��Q��7I�G|�c�[Ā�Z��:e!����-5���k�c yA����:m��E:'��PBͿSd�,�f��2[��[��+c��ǵE�t���|�,���]��<p�]��`�j�,4%�6U�U�]=���zA<q3c�����$zt � �=5u�m>1�Y�ŢIB��#���\ș��Hc���բ!c��=0n7�����yY?Uo�ܗ�©pi��1E'�S}A
����F��I&hᆧ�w�4y�N��?� ��@L�<	��b��k*�D2b@�@��K�v�K~5ʨϪ�n+�ȭ)-t��I�
Q.F�?��ԁ�'��S��{�����{8Ĺ6�5�u=�/�eŞI�~p���NV,?�!�*����(��*�@Z���o�=���5~��_M�a@o�O�l�P�/%s�����&1|�9�z���Ʀ����u��v�"�� �u��d#��u��uD���%�^&�X:��O�bǜ��+.��i}�L.�P��\1���`?@�J��!$��k��YI�2�y￠���/7~`Qzh���l��-4�|�O��L�
��8�m� 9�rbפ�?�h�0��4����P�*G)Q��A&[���l���A����G�8���K6^�OwAe�b���'�^a���5�	��Α�`|<��R�e\c�Kwww4y_&� �+�X�sI�}s\���R㷽�33Y�ܽӺ7�8� �m��M�{�<�W�C��q[�ӏ{ �r���o'�?(6&f��!X����Y��.�sC�f ��k�#	��Ho���z��q��H��4avg�N�5������7�BO'�F�?2S��ߖ'���<u��� ���%���2��+�ٟ�r�bD������J�Dd��B>Y����։!��l � ������'2�cVF�,}-`"�=����F�[�O$�%6~|E|v���%g i����@��x�j hh�L7EӴɺ�?455��9�v��/o�}N�Sk��^Ώٱ�������	����RX�U���3Q���Ca�ӹ]�Ļ�>�؜���C��"@y �a~˛�����/ ��i�/�h�,6�>V�S�Ա	��3�ѥȧ�-8�����u�͈�������«{���T��scC0�y���jQ��+K������I���6x��Q?.c�wsž��e��B�� �Ţ��1l�)]%�����'�[:vj��U��c�:���չ������y���D�{��x�	:��zbќ>,@��������%�]��y$̼oC���Q�@s���{�D,GJ��_ю�UZ{������7o��y��ߧ��@�E�n�/���y�~����Q��d<���}��&ngiɫ?���HW�[&2ob��-8/A�FC	9X2k?)��>�����1�x46��������s�/�p�����'� R�m$����/$I�Ѱ�N�	���M|qR�_-'�u2�L%������/�1 �\_�s ������9�\]TTQ�iii���!$$iiP�c萖)%AZZ����v@��n���|���Yo��{��g����qG�G���L�A��������h����������U��Ȗ�C[�~�����Lw	i�i>O9<6Pw��qh�@q�{�ݸ���}#@��3�5��;`x���,,xy"�̿h�`��ź�M�����Z�1 ��W=�����PǺ�<�9"�6F�9]�f���a&
a�o^6�l�&�f����<�8���oj�ނ�y�T=�I�U@�^,����_�)p��PB���]rSC u�G��o�k��Q���/8,-<���e��kN��9ͥ�߆������		,���ee�'�o�Q�DbO�K�N�8U�"�(x'��%	,�y(��	�k����`��A��V��cj�)E���(ތ�t�E�l�z�������ټv-ۄ�)J^t� C�Ϲ6�����x�G���
��2,=G`S�8��#x^��N���i3X�Р�30<c(��r�_�o�ʠs�i�S�-�r?�*h���s���B<�s��گ�fi�֫œ��-{�(�	�r�4@�e#@���:�D���q7�e��9�{�Ü?ȅ�$h��M#��Yl��\��|�����uY����`���7�R<֚������e�cp�΋�ПEL� Ӯ�]���!�/<�%����޼�3���	Qo7�8���`����/��H"@<_w������8��cr�0�<��k���i�y������V�<LqV�����i�O��O��UP����lf���D����F긲��Y^_]�������G���Q%w���ݪT=�3�����j�s��d�?��;P���0��o �pD�KK��(�nRRR����ro�����sj��f�e����y0`�4�V-�c�θ�s�`6[r�s�~U�\�S0Lc�t���M�I���`�V:���$�yG$�-؎��J]����y%��ߏ?�Cޔ�������z�O���|����ޖ$u��Sh�߬���[���=��i�[C̆R!G]�u�5�來��uh��9����߶�i�8%D>���P�~K���r�����u|�~�f�:�e���˵�)��F�32Z�@�����'�1�&��EDDd- kn��3!?��1����:�\��_$�IWfb0�I#e�%��E��cIW�N�!xX� h?���/|����؇Q���d�������5b�R?N�rѧ3���={�+++fs��"�Si.���(:$�qG[����;f�s�� \�ZG�h�앞h�m+Y�A�U�$(����j�w�����Jv��_�@0q��@�����{e澏E��੏ߥA�a銅�e #��c�D"<����7i��,�Q��#0��x�\���ô����C#��,�tu������`S(�X\�(��S@��t
�owt�Y��7+Z8��x+ ��:s:!��ju|ŋ�]���. ] �6a��Ŭ�w�k�<���!~7o��r����3<��O��>J j����\HS�R �&��è��]2e�z>���hF���� -p�*Y�hc+ ��P2V\u��̜C��s��" ;U��lRB�����ّ�0�{���E���;�������������#�7)@�6���M����yͧ��/��};�N=��`:�I�
?8�G���3Z>qU�C�j�x�$�e����D�@�>���#����9�}�,���u-�/DA��k��Z��2/�r�[�b��`�Pfg�-��3�������e,���|�ja�����+�v�H�� 4��Z, ��[�s"����_�>6�ڢ��6�:圣�в'��=���T��v~~WN�_��\H0�
S��M;]����ͷ�`kە�ƧMIM=�-IШ����r�9�fd̑.�{F�Ps����O�ʂ6X�R�c1-���8���d+�OTU$�����;�W�q��y�(Εo�Vˆ�ّ�����J��>!��As��l�������� ���'a�5�9��'�qL_J�a<�$XE�+񱀠�ua��/�����V�sͭAQy0�\v�ӑ��._��liGM׌=�M{�7��8������\z^�� ���@c��hn�6�a��ܯ?ò1]/k���Cw�Z3��Fi_��x��x� #���/�P(��t9�� N� N#~rw)@�
m`]�8��׮�`��А(>rF@����������!��6j3�/?����f6Ld���@�&3�����fYIc�CL���2��
�	(�U8>��-7�����=��J3��k1�l�eE��2�!m�$��:m���.Q�����K>4�D�>�|�NƏ�E�x	=[G��l r�͠���g��to�@�5���|V¥���YE��V����J%s2�%ș0�����b�6d��=_����"|L�|ߘ�B"�N���<���g
�?6�����1�����7o��?۪�4۷!�a�ͦMs� �md�M��;����a�m�	�ww?�5��Z�7U��q?�Ā9/�$��9�5���_]+����+�.*�־n8���&G��[I{I��0D�̓�@Pz�k����]k4�	�~w�ԯ�W��>E�Y��?��y�����g�̠p��`����AN�|KS�fL+3���ȐE��ŪT�f�^��3���M�ZػE!�t�%'"�r���	P!Q�+iѡ��������kP��b�
:7�K�<�r�Wk}�x�"�>Ǜ!�$ }	�cB����e�Aˌ
Y<8���mԾ��gQ �e���@Ҭ��|��!��汽�6��`1�ʢ���c����tO�C_eY_ ���/���UZ���v�r� ��od����!�,BZ�w��_�4Bi]{a�QI����l����V��Ӓ:Ɇ���;[�,B1!8B1�@��
L&i�V�5�~yq�]?��Q�i|� �*�5W�5W�d�=���닧�?6�	�s����-�z��:�Am����>�S��(m�$?`�H�����b4�� ��R�e�@�y.!|O�fLP+�U�^��5?���t����:�	�%�Ķ��א9_�9߫�^3�A	j��+ε���(B���dU ��Gz�	��6[�">����0����Q���5Y+��Ţ�4��,l<En��<���,�2f].�Q:9��5�R�n�u�����GZV�#0M�E�+�(˿7��=�T���OU0΍��,�vu�	FPA� �pw���6��/.����ĩ� �����e/�
b$H�G��"��b��#�,Mܜ�}���:�����W����:��)��C���BB�H�Ж<�l���2�*��f=��.�@%��S}��}���o�Ɵ3�K ���6_7��2)d��e�W�2�	���?�H�9�۰r����o�r��8�(<�ZZZ H���l��Pv�j��l�c8Ŕ��:.L$r�{ �{���n�������Tb]U�Uԕp�dR��d��d8�������g�����X�5���l7G���Oۮ�^����bY�vr�9���#jdr ���0ό�'��vbds�]i��r�)`)�~��g�"��
�H�[�f��.�Ӷ�Ӷ� �j�l�}�C�k�7o[�ڜ������>��ZKꞩ��C\{��uA^��\��;��0N�ȣ���H�@Qx:�Y��!rc�M���b�朆s�bHz�A�C?TL�
y��.j����̊���)���s��f����s�@��8R'ͨJ���@H�� �{$6��Z�o��_�@��?z��Lu���ņ�:�kO�M�����KV<�'!)99�1�UW��\o譱�ɯ�.ɸ�	|�q���k.~*I0���K���,-��+y�\�O(��U���޷o�ހ9�6��%�.5�?��j $V��T�3�333�G�Qc��+�	~	nzA�����ypZ�pNs���d����y���P���"pؐtk�BCC��ۋE#��#��&&&v��"_K�MOp��A�OO�1x��y3��𓷮���u�x{���m@B	U������z/^䲭�	C2&�899�~��N܍�JLL,稡4���$�4;1'4-"��w|s�Di�}�V`����O%�m��_ǝ�JЦ;�s� �M/�"�ܓ��C�꣎�9���=ۿ�a��c��"��"�6�����t�$��h�L�9SGī�;�$F���)�ÎοA�������9c�1&���hS�o�P�>��"�5��*cO��G��B�'Y�<�B�=�j��sr-;c�K/�Rv��7�ɪ�d�ڏw:tj&�s�޽������m�����@�pr�X�� C|��x�C���A�ANs9F��J%�x+��f3�Nj�}Ԩ���1E�H8i�'���>�H��1-��y�$$����f�uϽ^�h��#���Pbq����y4���bc3�=�J�yxi�#�ڄ �i��6����zg�=�E��d�����W0�V<]��ASLz��~ERRqO��3=�r�J^�/էn+;�>�>1B]�o��#�f�b���#"n!�8�z	����hA�������gܓ��՝�Sl���7�9M79�uZǚi���X�S�7(�8�aȻ%ZEk�h���`�/���ʒ�$W��r�c8m�:�	y�r��=�.���}�G�T�+O�9���s�o��X������"�Ⳙ����+�ׄ�Łdb⑱������(B��fS̀���)���'�7�o������o�7��f���ntɕ�6�?<\���׎�~w��Ń� "D���i�zm��$b콘7�%��	��?!X���G��39q!=��9D�R��*��6�&���7��aT=2mԫzĲ��0*����s�J�� )�h�Ua�lz�bQ檅�1y��i�N�;�̔����U�.'�±l�*�&n'M�m�ZU�T�o�%��G��o��~�ج��߁r�g�O��Wh�����I��E�O�D����^|PKL<�n9�����jy�E}�Ӝ��Դ#6æ?	��8�����Z���܈��Ҩ�H�?EWg'����WH1�P�;���X�>��b���H�4}�xv�5�&y��o ��g�S0�C\(�9�zO{TP��р���")�sS'�rw|Í8Rv��Ɲ5�k+%WR����AG��j׵m��bK�~ttD��Z1����f(��e����q���[��*9�	�2	DjFo��8��	d|c�P0d���GY<���c�S;��\�,�j���GO��ku�娍��K��M@���	�#��ǚ���,�q��x��^j��i.�0�{Q�%=���V��J"k�����k�e���ݖ�p�2$Ff�ǝuՃ��Ez��=�;N]Ӎk�I8�$:�#Cj�b�0�T ,��l���𚯽���g9XM���Ǆ|���qky�xrZ���z
���SZI� �zpk�\6�����*���������3�MH�Y:���b��~�q �t�G
�g�sV��b�����bVE3:5��3��q��osoT ��?fSc%~R�����&��?y`�W��KY	��'���`��:�/�ih@�0dƒ*�q@�=��x���Ա�1��7g���C��4r�ȇ������r5x$�f�b��I.�*�qb;��h|�������NR�s�s]�{�%?��i�M4.L���>�][q���늌���u?���AoS�`�}��ڞ�Ƞ쵑�Ww.|p���o>k�80��p%KW��66Tg�����}! �z���_���d��5o0�fг��E��^@�����l簇4|)�G6��\��BZK����D����AxSȒ�n �;1���MT�c_欒��%�����B�Q�����X�V��;x �{�L��\�a��#(J���Yb%��@R�!�u�L�WjA>���.��$��<||�'u�+�����~	�(r2���T�lEV�n�k?;��C�&�����6u��לo
��\k��EG[Y���q���(?����9j!��#������0%f�~:�D��) �bo�>**d��G�
���t�fO�r5��h���q����_�5ߏ̅/�>��U>�4��
&03�y(s	���Ƹ���[��1=�O��^�_���yPݽ{7P% �F���u���ݛ���&����&
#=�L!=񌰬Ť�bsNV����&�>�K�Q�X���q�ˈ� �;o,>^l����%�jf	��F�}����-Z]�������Ӵ�^`�*��4Mo�.�m�uD�B�6����j+�X�*/C-'}�X_g�,�_n�� 1D�@0�Fyq�ؘ�g"��q��u| C(�?�ќa�o��X��1� ��q�tCL�U�����^�b!N��4��de�pV}��>I�(��fDq����7���ap�Av�zɤ0�E�T}ןfC�:b�½R�mI�\�3�A{o���N��wNfpÞ�|�K
&W1����ff�Mlإ�6=�K�|�����Њ��C)�襵���n`�bf�sc��0u��T[�j8C\/���aI�K�I7�Jݹ�B����[ElGw��g(Y�4K��K���h#��/]��/�5�z�z泙�Fnj�i�
�f��A������X��PX��8g/,?]�P�V�0l�xKCd��0y뛛K��ܷ%Tr�Oz.�)��t��Y��O�DOK}�է	)ٖ��b߮R� U� �5����)�=�AE�b0iB���`����	~��Z�G�j�F�ys��j�ʹ#�Ps�u%��]�n��e.����1i^m�25;�h��==�P���R�W_�f�"(���_@�X���O�ZK*,'Q��\t�[�wA�{��-�J��=K
1-7��[��U�83�X�����z\�}r�;Mg�äG�[&옷y�h$�.����NOV� Z�2d:h�z���u�����wX�r�v�j�{���
�IB���XVR�&�.��h�s���ޕ�a7�O�J��u�I
�b�zf���;^�]�zA���~��6Uz����v�vc���[C�=`z11�>>T2�{���lJ&�u������|w��#�a�l�g�q��,T�	L���p�><W%�	s\�]o��'Q�����eɺ��x�����$Z�ӝ��?�9@�>W�V�W�6��2iE��մ�����42<'�yy��������r��KN�
ƭ������z��^�L��.�"�ڵ��:���J	
'��d�S$�}��J	��s����!|�djk5�����T�ٝ� Ȭ�A��6'*��^H�;�̥�����1��܇L����3�qo��8>>	?����{S�"G5�������aītL/������*ʞ�V��@�r�.�@���mZ��ŝ�O��v��7ߓ��88�h`Eȴ'���R8&P������W�#+����.T7�M[E�0�DEp�����G��Y�N���v�"Za!�V���X����#��>$QBw*�av� �)��y�7��s��§��oWgˌ��eG��0���5��'��)��K���<�+��$�RL�H�؞gC�Ƌ�� �:8`� z`b2|�6�8����?4,
���p�ܳZ����|�r�.Y?4��9��;��T�~ػ��l�x�Wb�ԇ'�@��)�PCC5�Ǐi;8���PeՄ�^Z��TVWW_���L"jͨӴ<V�-�2��G����@�g�B\P�~���Ҙa��
l��Pt����y��$V���VzF0�I7joooА���og�Lh+�R�,�^󞪞�Q���J	��u�=@	"�����c//���Q_ᲜBv999c�P��c�����;��##���CM�Ӈ��_;A�,���:XlE�5biF�9&}&+�ǄhQ�]��	QdՌ���j;iE��S��F��[�˪Qtm��PS�%QS��VW�_IEEJ-!�%�B�~Z�]�Pjl���.�c#O��!����X��@���ЮP��8�[���l��(*|e��!\���1��'�>Pm`\VW-���\'�&���-�!���FN���\`�Pĺ*%Ov&�d��p���R$���۷�_��x�ܟӞ/�K��a��啕�5DH7՜_S{ڜY��}=���2�r�̯!�޳=�7{Q��j�l�V��-������l)�,A6�s��=��a0�V4.z:M�c�D 	������j��NJDD��XN�,�����M��\t�푑FA�DFLD�VP6�Uh��������;�h�>Ph|�y�����V3m+��nD�v���Ֆ��Z��ة��Ï��g5�[O��(���	b{>XQ@������yH���t�Aۧ�>��)4!�#_��x�EdA�Px�� �򲲀����X��ZIuM�=�Fޓ��6=�v�����mm����脑]�&s�a�N��<8( ����r���K��K%B��'�v�D3��˯�G.=<�<�p�[��a �g�^�U�s}�����ϯ_� ���/����������>��V����b�������[W�q�C���`��Ai-�(=?eݢyN�,ݖ�4�A��|<m��{����^"H�-=�V�>޲�t� �Ǆ�<������9�(}�#u?�a���)�a2�8�``KƳ�m����9������r';�}cb$��+�.%so����6��g�XX�����0U	榏}s�W�s]D#�aQv�W��{g˯Tn���c��efc&���!=��m kB��1 U�!�<�P�Q뼌U�_��C4��N���б���ۂ��o�o��k�P������4Y��%� ��,9��I�no��}���"�v*p�؉*��{�)��)]��S����ыB�:�P����G�*kj�uc�W5狐g���}L�'sz�XF�Q�@*1��i���{�.j����ۛ���������-�x��}d�y���M�\h��))�}7B�����U�i���x�E4��Ď�gn u�)c{x���6�`6����#���Ij�^q�;�١V�dySS�֖c�'����vI=VF�����qv~��W�2(��s��őZBs�Jkv_{?eQ�2f�=�g��f9�|����|�O��C:I��g2@� �\��>-'�ӢNQm���@?lⲴa$J�=�e�UG�S�$��N�ՠ (��"rPia~͉��$�iRSSuttZAx�s.0�l�?��%]�j����P��,/��,L�.;�>�x����Pe���[T�".�'`�In˝�E�hQGQ���^y�O�@��Ү{t���>�IIIy<X~��*c�A�=�����z��[�ĥ�E*�b�%H����L���}g�ݻ���)y
l.&RA9]a����u;��N��Ha�c��pC�L$ 7
�\+�t��7�
���Z� 
�İ���tB�p`���Tylr{d�}�P��$���O�WG�L���^eCNK�"U��8Ϫ�)D�	���n�?�=7/�UJ^�M�o��q�!Ҧ�mp�)G�k�?��#�mB�#^��	whl�ԗ\����8[�I��Z��oc�s�ޭ(?#5�,�%��w։��:��Y�X����i��<��h�Ҥ[zl g�u�m��*��l�U��_x��Z;�J��`�g�Q��]-y��hQ� �����%lz��.��yr�����d�˳Ci����]KK��:��K	�c{{�����ӛ1��ļIɸ}�4�{LOyJu�s�_�v�N��܈�&1*�{����ŵ�?\���]J�t����k���MvU�.����ۣҖ�[WQ8��|8�� ��:�!s��*B`��\079%����1^�P��
�0j|�RB)���Ŵ`ç�LEl���)��]�,mȰ�܉��΁3�VA�,�'��q*yb_�
�먺�=6��Gw4� ޡ6�k�>�o:/4&�h�R�ۯx˪�HH��3��j�ijj���ε2����i<�{aa�׊�olj��ͳ���)�x�<��BZ򱾓��>)F bґ��<�3C���TVYtO�X�u��,wMMʮ)�O��Q�-SB��uY_���z%�ax�X��dn��fd�ό�X%����4�����h<ӊba�vg�!k�m[�_51e�ñ����iwGZs  �ˀ�b{^�P���,�@n�Ӂg&��c

٧��µJoK��^���*�����·��Z9k�����'���|T��	?=��/|�#>7�`Y///oo>_ �o�^��#�+���H�YOo��C~lQiH����v�2��+1j���ڒ~`q[
!<�޽L���k��x�O�UVVacr����^��6S����R{}u��JC�X�7�w�4�\��!,}�Y/��J�О���&%��"�e��2�2�6f{mb��e��O�J�X����+g·rZ$:n�\4�;�G�k�K
ll�Hѣf���+����7����1P�%�IKK.,,�KM�.���!6&(�6 m���4�ޫ��
G����Z`��2�d�D��d��ɠꤻ�a�*=β���B�dJRuE�<�����v�4�f���R�B1A^M�f	cl0)E�Dk�ǰ��������A<�FwA*�Q!����+�1��hX7�DX:n��ߖ� �%�Us ��<�ܼD~��c�G
�Q`$/���Td�]}��w�!�%N��־xZ7���s�����r�� �a��O
5؁�y��ϊ���[�!��Y�C�޽��֤������~�����p������ϰ8%fߨm�bC�`!�Mr�Q��_t@,�Y�t�!��o�W����j����b�ԭE�|s:��
:��/�H���~���C�]��Ԥ~}M(�-�ua�a�aG��������� Qq��%�	�5�ITc@��ת��|rX��V��%�V��V6{�~��gQ�dhxᡛ�WL*����)��b�w:w����C;�"B}7F��n��Ο�u',t6���� ����ƼM�r�O������:"�S�;�+=��U����z̢�{T}愇^�k�g�;p8��� fww;��lm9,�O��*�ģZ�s�;%���x���t���	�����5���t���w�����G7���j�I_�	:���")�o��~�	���F= ��?��d��C�^}�a�r j�o�r���UO`�7j���.S��u�������̥�����QU��ڍ�Yd�>�-.�����t�ֳ����N-��c�g#�L����(�L��{V��ɍZǟȀ-~�\m�#�Wp�V�v���@JF�S�9<Z8���m���ލ~��g���kv�CC!��R$n�s�@��~$<H�=��g{H�t�)�����gN�߮,tI)�F����f眨���H���x6l�'VZ-! ��>%mB�D�����U˳,$S� �WμΡ@@ɐ�o%��S-�x�-H�wx�)ܽ]�����hl|��S�m�������b�G2+���d}6�ͭ�׊�F�XY�e�Z�oX���;f�8�����xq�:j���bo�thyA/��+u��bn��i����9Vz��?ML��ߋEjz�d/���!T.��j;��n=*B�ݿ?:r����r2�)��,B�NE�s]U����w��#�s�qx����;e��W�E��Ck�<�ct�έ��_2a1f��|�siT9o�0��P�*�h��e��H��9m�YW����VVV���a���Y�xAܺ�m?~0ʏ�[�ŸG4m���O>�D�}`�r58�|��,cWױJ�����D�R��Hyt�M���������3���:j�����T5.�3��.)|ۨ@�����ϟa���3���ʣ���m�<���pV��[F�z�&�5]cx�W��mU o����3�!䘸�(/>^���<)'8Dl��E����	]:G}����C�佅HnS3���w��2P~kkkra��ώ
�b���������c33JJ�@�:k�Q��E�!����������+T�닼�B�_��[�n>a��c\��A���0u~�Y�moG�����_Mےr�\�UWW�/ܧλWS��+Yw�?�v� 6������<��깿�xR�՘G�����#��m%6n����\�+[Ĝ�;K7�S"��ڞ����Bl$ka�#��8�!�kQ�:�@��*�$�Y�oͰ/ ;666i�)W�����~�计y��+�W֛�oƖ��7UmT[Y��^(	���ӡaO�T>�W�
��k}IX����pw3�DŪ�IP��>w��+�Y��4��<�HJ�a[N��fK�g�ߣ�2ݠ�3|P�p)�n�	��3��Үa��`A�|̷>�.tF���n�GV�,5,����.ZS+���"���� }g~�+��hhp���>��&�g9�����ŋܭ��?7�+=�r��p%��ڵ7l9��I�3/����K�����z�"����nwh� @�):��EX��%��Ǐɩ��J���\Vt�q�r���A�xlD�Č�r��Ub����vz����~_ȕ}і2s����)ޮa`Ca�N��.�����LS�u�WY�{܁N45�������L���|u��/N<~��=� �o�*1��0�g�������1J�a�}N�+�����Z��L�\�����<���c�t�9�th�q�E�2��84�#� :����Ʒ��:���bc�LL~��x�͉�ɚ�H�j�*#᭏�M��8�~ό�{���Q:������ַ�]Kd5�H�k��m/E��!�6����TR"�3����Ǔu�"���]�EН?��B,�V���)�����p���afn��k�NNx���<#��ꃄB�G��Hm��
�m�G�Q��0�o�a)��q~�1q�w�*_�f�/;;;Z���˕|�dgss3�(ub��}e0}�m�*?�ۊ�Lf��q����7���C�����2<��Hs$���?h�U7��]p=J[/OW2��zC)q?�q��+���	��{�: �����\]�q�j�^)l��@1"��{���H�JϮa��BT�����"+&��S���[~9그w��k:��o��ю=�{jht���:1���^K�9��6�YD��A��N�e�_��3���J��QJarpq���~�j�<��@�ĵCs�z-Fx�b��KQ��R���ݦ���f���1A�n�BO�κ�Co5j�_��G�F��Q2vm��+F!#*c�����²���uŘ##�~��+�e�H�8���'z��Rq@�O��A{biR�j�(-��w�+mD6��*�����5�հ�rc3���5Åm���=�I���������jh�����5o	=)�����,����S�zAY�Z��Vh��666�"}#�B�����ۗ�N��<!@�@?,92�z�A9A�2�e��w��ú�m�]Xr�0?n��PQ�l��?��& ��!nwӂ�y��JRq	hQ�\���к�7�J}�ț�����N�=��1q9\�l���q��K`Ao�c0��g��3|v����ֶ����_9(�cg*Ǵ|�\�,N�YR���a0rI�S&�%��;��@E¨��-F�����c	IrZ�V�'��ޱ��dK L��̡<J-��3c0��tk<�nc7W���\V[ۻAr��D5U��%�H�t~'40:7
�JX�NF�
Q�����@l�'��YQ�|�za�(��hl2��[��sx{b��1*b{�kk��m��'j�TǢ�F�Vp��Э�p���[����;�##.u�r2#y�6���|0A���󹠕���t���C]�{����GU�r�l�?)#�S�fKT�kh�
-,�2$���~�����Z�K/�%2Ad��y�Y
3@QbH-�Ņ�d×%H�G�:_*@�O������:���]5bw��'u���-QJ̣δ��o���$�l�I�M @�F�F���۔����+��2 6<�]���ſ?Ӊ\�e��[�	����5s+�p���H��Jo��Q�����]�ä�_!>��?���`�%�@�`ra	�8�������Z���3)9�3:�<���,�\Ge��m����-x��<���`��ҼHyAM�3����N�x�^de�]@��	+�NNI�qq������;�(�|V��XvϷ
�-��2������ �����Ez�vPw��PK���3�FZg�Ұ!B�/}F~~J�%X�y�*�*v8�!�b�H)��_΁=m;�.�UV�:_l���X2�~�����VC,���/ ��3y�����Cw��w�{뺊|U��b���]��
l�uu�s>�v?�679�{z��Q٘�zھ}S��r��R�6�cE�v�iO����>,'=�u[S�:,ӌ~~v楡x:G�9#����K��}�?�L��v]����H&T&y������J�E��j?���-�u�tC�t�?����e��vi"nX�Mκ��V1�?�?"T 1���<0�(�q�U��M�ZO��li[6�^�JT�����q�fA���]e�<����#�_�8̤�$ݰ>���h��qnn����b����R�0ȧ�_�04gd�s��D�V�y:��m�с�����Pw�`����?���ܱ�IS`�C-���'V�t�m�onn��y�����F��������
�z�NrU�9ץ�P���Δl�<a%�ێ�g|��������.���(� �n�I#v\i??'��9ꡮU'F���/��Ԝ.(����5\�9ȫ�k��d����#�hq�pϡ�=� ��㈭`�J**^��7-ƭÉJ�H�h�>�#�A�u�EA�9ߜ3��y�2�۾�7��ν��HQ%�L�@�]Z/:��p� FV�cf����]o� ���0Ă-J�cY��}�8�:ګ)XƹAI�+ǹ�eW��{�����u�=,z~U��#}��_S�o߭S̽�ҝO~(�,A�a��u9�~ǫ_y'=���Z�Ft'N��{�����mNH�O��x��>�P��p��]�F{w7�u��A��/2ׇYg�*�u'�ж$aS���{�4�.�>ȵ2uv&5������|��i�3`�#l��k@36-''��OIej���XN�ښ�G��qy8	�i��tli�;����s�p/��_o��kkV����Z��t~�Flcj̜<���v�1������X�єGE�q?�h R�K˧��C�orQ*�[C�R��jHxx�������c�W}6HI����� �A\~*
v�p��Z��xO��������_͎�bz g�1O6�
�b�He4�����A<���\J �ы�Rǌ����y ՗dk!6��C�Hr��m�u�L�0 �_��ƭIBMZ+8��(�B#��65E�Q?�5���5�mJ�u��~�y���o�! ��V����z�[�jB<JK�%��{�n��4!o�9�"��VA�\[s����
,�~��&�{pi��$,7�ϛ\�Ԟ:
N �YW��+F��~���p���87~Yu��^v�3::*-h8�T��%�׆p�	y���2�Ԭ�|��q�VJ��H;ͪ�qZ;��W�-ש-�G㙋�����C:"(����\oLLLo��9%@2���n��h��Rq�"��ߋP� ����9a`����%��?�wl�?$�'�����O������ڡ�;P��F9�b岁�"/,�ʵ \*�
��n��>k�ӫt��\�"�f[â���g�v���3�''B�2t�u�ǆ��=�����Z����[�a��������š_��3$�*BI#M�����瓞?؟�^�\_rl@Cub_szYwy)�١�˕#�O���+?� @ �b�:��s�}��0;x�\��9�4�f#�Uj�4���Z��
�֡6��A���]��OĠ%�}��t����L�C���2U��S�G�:q��_��,Yp��y �����{�i�F��L�/��܉�1h�$J�2h�th�%( ����B*��R�ƞN7���@Ø\n�ڪq�*���FE�)�C/�y"��3�J�Q��N�cl�-~beo�@�ϵ��B�aRj�&�c_B����{�����_�	o))+��85$ JDA�G��5K�Kz�0�~jn���x,���u�q�ş�Ks�����F�$Uz���葹Vͪ)��(�d�9�<2Nr���IvI-�#h ���(�)��_��QFm�u <�����;���|�t
R\��u��U��X���:��r¸<��#����j8l��9��ښ\@�$*�l,Z���:߉�Lׁ-`��~@i�M�����<���\W�Pr`�:{��n9wNpa!���n�4��#�x�"d�-BA-���~��;N���YU�6ŀ���a����q�'��3�#�����"�|/}�iK/u�dJ"�P6��
;JO��l�RA�6���lL�N�/;�n��X��KM\k�!��'��P씦o[��n��X˘@��XJ�S�T�09W󢢢���.�c�NU����m�?�0�닒��Q��q�-�ؿU|]^QA��P-q����:q˴_����5�Hkj�n5^�Y�ت��U��<�¨�í��{������(�ȩ�v����}��=�-�A}l��E���O�Z1�l��p�z����=Mt!p�v�f��=٘�E�B�����Zh-���	�V+�x��`u���'�.���T�<��nw�� ���*�O��t�:Q�E~����=������q3�.�h����{}�U��Ü�Q�A��Q-�[t��a"ژ{P?�B q�X�)`�b�3��>,�N1� �������A�o}�6u��5�\\R��O��;x(�.�:���6�
���~����1XM`�9��<�L�
t��Rt��n����R�z���]��.�uUJ銱���<�ޯT��g8��ed8lBY�ϯӗc��,�	.�@9<8���`'1�c^�X3<�L�HOϢr�S7��M���H3K��˦��F��$Q)҅au�W���f�*��oo� �d���_�0��{�ڑa��v�-��w "ם��t������ro����ʁ�bCH�$G [N���=.���ˁ��ǶZ����Z�4c�݂^ �PQ��}}�?6 �ĝ��v��Z�` �o� �\l)�"�����nnoW�Xxzzf:�U��D��ޯ1)�(9�������( z"d���&�qC���{ѥ��N��P��!#�ƶ^nnn��跱G�t�[�N�WzC�rt��2��v�<�ꅅq�I]�����T�5f�u�/��B�F�v�8��zq~�C�S�����~��O*E�3+��d�:����d���,��JV�&�X9Y!'����3��N�O����ݺ����^���?���y]�4gD$�S�S���;5/��!U�P��_���G�����tx/��Û��撒L��f�3!^Iu����w������1R�we3��L�����t�޸n
���t�ni�MMςQ�s�#S�U�U�
�B���S��7�9���"� ��#1�&&��7g�eˀ�9�iSg[�or�x4�]bΰ��]�\���_A63p���(=h����@~oTK�Ω��K�A����RWQ�ܳAI�5#���}�U?�G��0�ozr%���-%�ס���h�V/i�'�H@4�r�O�n���W�~ax(8��vm�e��{��!�䝝]��r�{�V~��s��!����N�- &��k!/>��(��#i�;Zzx�PSS?�oΘz������ڍ�0Y���(����^oc�,/�c-�$if�M~���9���I��O��)wo4�D�oXC�\<[�Si�ʒ�֣���L���ZYM�t��?�:5�(U��ca�~L�ߊuV���F�%������N�M3���&E���Ӟ�w��M{�����N2.�����ߵ�T�5��{B�r��51�X,��e�>+"{�4hnk[�"��SU[;�����fu$c��}�x�V7��,&tN����}~�jdÉ�[DW��r�,z*?q}Vm����"O�I=������r�E�jz��$��2�|�ϲ�T��p���NxW��e�����{2���z�\P�}�'#g��F�᪥��uJu�"U�7V�p�5��!��m��c���y�s������g�(�g�w���ش��N����̛�j���S��;������D������=��ߩ���'#x�����_}݁۷e�w����߷�rpϮ��G�9�t��,�\Cg9&�a��)�(�:��Pp�#h#�����
�,�TG���H~zT�U�f���c"�^i
JL�q����WyDI��3m�<�H����L	E1w�S��:���/[����kr�k�㔏NZ:������R׈�c�7��<���S��y�������V��n�3G�ܤZqb��㺝z-��?oƺ���T#�[�++ww�A60�
k����R��)�||�=/M�3����ƾK�Z�j��j����m`�ٜ���]H��sG�6b
*-u��Z��s����� �-zއ��-?�w
�>�4y��ڈ�O�C\�r9&�>���Q(��2��ޜZS��F5 �8����Ē�h�ν�>����������M�8(�	}���d�=~��ǿ��&��(Z����Փ���j��j�W�v������J����V�#���KJ ���=�鴏���~6��G��B�:���O��y���H���w%� >l��=�W{�+@K�į3T�ҟ���7=Lޘ3���hrPE��+�3���,(QT!z��f�<l�[�t��aFx��!nr.���\�؅�1;��y�(�B����e+Dh�U�Sn�sƐ,�u,�l64y�gk�g6L��r����ʔZ
H_
�ٹŝ��/P�8S(;���Q\������!M(_��}���Y+�7t234\-�C$R�un�tM��pt�8(z�Y)�ˊ$�`��H5��c���pk�ҫ���]M�%ݷ�KJ��� ���(S����R`[��D�eQUIb�ҍ���֝��-�����:J����ܠ�O��гe���!=]ݠ�%������,�Å���9��FC��:���m��l��`0��YxCo0? 2톎~!%B�i�QK���q./��_x�6+�*4�V�YS��*wGXPJ�QvVf0�6/^�H�Wo��V�m׍W@�Z>����&ϥ�ZH*1��_��6�gA�j����שA�܍�Z�z��LL�~�l �O�T��+l�����GAn�����=d	�����4��gv�r���)]�]��}.d?f��ż�+� z�Z�4ٚ�k8!Q3�t�7Ai ���ŭ! K�.l�26��]�)=�����~���/�
%�����ᎉ�|č�e`H��ݿ�
刿���_��쎴��#���\*ְ�5�4)goo���Orp�[ A��Y:8��$ߑxB���wo�5��z�tbnF|SGG��j����#70��$��I��i�\_���x�v0����i��'K
/KVyMX"�kt��m\��~
����(�:���e���4EΚC�A��L�yp�>��h��Ɏ
��7�!J�I�ַ"~=�.���$�Fyj�8>f�,
o}Q����_��:r�I����x�-96��k$���!�=����g%k�����\�XN{�uC�����Ov]b�p��ۻ���*�n������'�"BB�O�ހ����XPX�lcc�_���,��$nnn>�n=$upt�ep����p'��=�4���xj*c��+�?�����~£r�99U�\��LZ
l4�y��9��v�������*��o'/��0�|4Œ�F�窪Pp1��Y�ć�H���؍����i��������%��v�F�?]�E���hV��X�$�ag�\��p
y���uA��0�n7�	#}�o��.2��z�7g���8���a�ܝ�e�f^2 xc�6�Q41$�2��u�Zyf�zw��%��?�r�@~�6��A�9����A���K�NWRĆ]�LLL���s�J�Z�#77���I���!��������-pj�G�1�(^����((�o`�D�$sA�}�9Ec�e36��E��>�NP��\!��ѩ;�s�m� P�M��vǲ������C�k�� X�F�`�Ι/j��oL8�W�z_=��NI��)h/xq��;7A�ip�SA&���+E ��:�]��f�MA�U5�x�ￖc���A#���l��[oYp�u�U��v�Ks�昲^Եl���<�k�Q��*�����dU�4��F��6`{�p�����z��-�	����IPQ�Z4H��Rn� �J-AZ���4�	�U�A/z9/��!*���.�f��k'f�$V:�w�M~.��3{`{�'*#��_MY_����/�S�2��� ��Q��!r�||<�Y�񦂳���k��|?cu�II��Ys�G�o�b^�j��$�g}�Ζ2Q9L2���҄���E�/���I�!�/��/gəc�#�����W�o)���!w7�7'~�U�LU����!��}t�f>�7��CѺF��}�4�7 #� b��7��b��o>��R9��䝠d� Z����[�5���,e���	e�h΍�P�ߠ�����3�q���a��~�ю<|��	˭��H ���"��䇜����#W��}$�urŷo���Z�q;CAtf'��;�C��N�T}��� ��{1HMI&�O��ё!"<^��2Z�,��~��t[���;���M({�u矷�C*��x�8;WZ'�@9B}�G|�	�6p�����͉�<���%�e:z�4�R�>a��y"I�u�=����VQU�=JpG6�]�6w�i�v�8oP��/�D�����l��͠�Ԡ�:4��E)A��F�Ϻ�q�:	��ng$5�>?�a�f��g�dj��ai:$��ګ����]O��$�o��PGlV���J���ºb����ƿ�P�6���׫jj�z�$�'��Z��L��t�NA��Ҁ�D��l쫑Bubݺ>C�ZǶ���HsO�t,@�Û�ސJ�]rn��q�ҿT��w]�l�H�o�vthq��y��L6� ������7c@�3�	Ys����H��0���&uiF9>��[��]=�`�+;�̾|���O�#[��dāMɀ��!�6���P>eD# !엨��/����o���#���dJЇ��$�/̪�I����Օ��a��(>����p�y#�F�3J���|�����m�ad@r�ZDO�]>��km ���SPP�Z�\�HM~'���D�܈�����5��W)^o�WQ�����eGeD��₸��B��{F�i���_JG��'��w���@�#|0|���3ߊ�;Gѳ�uŜf_%pс�q������P�`�\��TG���n�)=C�5E.�}����WvYοxߴ�XJ���M��=D4�k�e����eb��P��ۤoNMM���*��-��e���N0�q���h�D�@��-��M���h���t��W�C��y�@ڹco����tKp5U�78x�ĝ�6Ո�0I�OP�~�;�g�v��-��绫�7(.�O?{w�o�Q:V���8���n�0o��fhZ���l�ߴP�ֹ��@f�>W?�~���&Whe����3St�H������)"���K#��K��BZ�������L�U>4:�)��;֧�#O�8Y�jz@����Ɔ�8���:Z�!{>�[��/�����l-�E?$BX�
�1V�k��w�k
g	<��,(���,Ҿ��ujjjR5�Qᜁ��{{�� _z;�����#Hy�������/}_E�7"�g|��)��Q��B��������Ǝ�.	�-�'a�0��ܱ�Nf�_�J�*�J(fɫBf�AZiͼ�ͦ����xc����q��`u��[��X�ζ�M��%��FR�,�z't	����-��������A3���+s�+G��Q��M�#�uE�{�&_>mk��o.�3�m�d!#��o{�߿g��WA[�<�UmM:��I�e���s0������ ?�a(������ʊƁWXEN�#�n���6�d��D�3�|�������K��R��9�[s&܌,,�^�{���'B��=yr�+�V?{|�� ����|��n�ЗČ�{ŕ;^g�(�ت�w��!"��;f�j��McY��<^��'{'�
e�6��� �������7.h6��Vn�X;�} ��7�������BY���`�,����z��P	M����s*�F�����Vnኴ�{GE@$��G~��ʳ����!MI�ss;~�(���?y�����uq m�z�j8;^���-&
h��Ð�o��䯍�۩�@�J�ӄ�˚�/����^��_�~��ߎ"9㟪e��T�?�{�;�I@yK��t��CF�BMǭa�O曕��Q3��eƍ���@���Ly*w1����U4t�4��*+&������_�w�ڵ i�h��
�!�bm�v�A�۷�7<�}�Iك~�G�.59�zsQE�����âj*� ����-��?�nL�`���@5Ry��;�EZ�?�2�u��YϿR��7�������g
"l�����ޭ�y�y����y}�T��2e�wyk��L�=����Z~�*�;���6���+�ӎ�w�� (��h���T'�j��C>1qq����9i�gll�c���T�N��+u��)v��p�?SV'�q� �zJ�N���H��[�~L��w�����|���ΨM��'=-	 a�}̗���p8FѤ�d� �G~��I*ŬA�;Y�n;�����-J�y�A;ۿ;>|�H������n{�6��1��5�c�Ӿ<AK�A��h/��:����.[-X�Ŝh�L�hSS�ܤ�=}�S�{	!))���Ь�y�|��sĎ��C��t��E6,@��p2�V����O�^���)�����w�ϝ����HM��U�q�/��0܃��p����g�j�\�|3�c'k���9���O��	���S�B��K<���{��R��:Qέ���޵PJWf�2h�t������~)�_�q�H3[+ʉ/�{�,,,J�~C�/�T�[-X[7VW�˗�omU3фq�o��� �f�4�h�y���7�EPt�xmL��W�>�|,(��#'�g}�)� �羅��\��%4�P�Pͼ+�����`iv��_)~{t��ܥ��z�]Ev�`���MY�}�������}�I���k(�3#D@c��
.&'W��CZ���:ؙ��T^"�9�4{�|�����:S��=����\G|�qG�2jz����!�6֊����$<vvM�ܠ��p�����!�21�^�I�A3A��)2�V����Xη����!�t��#
~�`�ُ�e��}�2q7�b�E{���]��S�Վω/������%�QίE�QK�����/
���|7����N�6ݳ��饌#G����8ۯt���Zn��VH�}aho�O��7m��om�%��S��hMjg�r��Ѭ�����W:I��ލ<�:���@���IWU�E����#-i�s�^x���rF7��2ߏ���#��'���ăa��M�q1��#\�1�>6�"\�xp�D���#�!va,g�i�b�`�mg�U�z;v;�.���.�*}Օ�Έ#��0�����t�{mj�|��Haފ�D������F�F��'���@M�&b��O�u��3�~���hcs�_�q/yV��/k��w��[�k��>�ja�M���h1-t���bSssLi��pJ�Z��'{8Х������zgD��`�ðZ����Μp�$1�M_`��8�h(XQATt	B�Q�]MXb��ܦ�����r�ӯL�0����k�H�z��O���~��k��w� #�C�x�Z�����^��{����P���_�����������r�ƟE����t��=V4O�+�e����N[�n��F�-�Hl���E�jL����#��g�YG+�Q\?�ۊ�7�l�F�@س�������0N�%	0�[�h�,�Կ��w�G�Cr��ozOzv�#w1�m�z�&��~��]����x��ܘR���Q�S���ׁ/��e�ɒb�F�Pe�Qn�!7Ĺϴ�^w��H������^}d���h��l1��{��7"���+[Ϛ�jof��)��h\��zy[���I&eǛ�v�!��/Uu+��݀�d�����D�!��3*5�FՋn2��j�'����l����n?�����M���I.���nכ�w�6ؖwV���w?��r����~#r�Pj�I�5Dt�i��c~C=>Rp��JM�^��/��a\�W7c6�>����"-4��z���j1�|c��@i|ì���w[���U�mA����Ѓ��
�f��/�p=V�a�&�(���q� K����`eV�B�&�U*[�D�!'ߎ�ר�����Ύ���[�I9;5���_l�#$ߛb_g�K'�ښ>m9:����Z��E�tlT^�%wl#��ן�ՆA�dP�N��'��}U:�aJm4 �O&�־Ξ�7�ė��)��>wR���8�49\�U*�V�-��p\3���aG�eA��-5���8i��������^��T<K����4| ���6�c���U\w���2�X�Ʒc�|��;2]�ğQ�F���wo�3��f�g:��D��)�P��=WItH$�I? Ĥ�\��fߥ�O"Eoͪ��z	��G8�K�\eY���[�. �n9��znũ�A�;?{��U�n%��\�_��A��fi)�(t^iY�/���l�<P�%�����B�++�_�z����ꍏ״�T�����_�%�t���o��pnk+�zf��$P�XB�Kgɲ���J=6�8����\���`��ܭ��;0Y=!�����Q�E���6,�J?�O�'��|M۠���T����9s�.��G� vTN��[���,���)x��W�5K<v#�	�^/����o� �^ZI#������.\l�<l��<Q��E�	�@ի�?д�[H�y��ړ�(u?���ޗ��/���Y��v�QX�A0�o�B��4=�_�-�}�~��鹒r�鹋�K�Z��v��ho�b]�%I�Q���(�r���9v�e��	[1�%O�Zt#�{�4��B�f^�'��oCNk���@|5|S�O�dAU�B}�����m�f���_��0%����1����_ט���I�ֈ��v�BQ��]� U��`��_��K�/��T�y������=:IG����y%�
�h<�399�cb�wp�=��wj������@|����:ڞ� )�mjjvU����q����@�efff��(3��Z�@�J˞�)f�;ڢ�΂j��߸U��q�k�W	���r�ڿ��=\��+K����� 66��yFHC�Z������WA�l�1��m����/�0���naE�c:�w|x����+&�Z�+��7{�Nq��+BS&���׹� �9Y�0�I?�|�R%�����P=1��-�[��~��2 �Gn�pw�$X��J��I�ʮ��O�I~i �>\�j�<�a�6a�U�F+Xwv�g��d���_'rꑲ��/�Mwz��; @�[YЕ�����r�ϝg1�?���tr�6�h@'Ѐ��ۚA{c2܍��Z�'��}y;W���/�� 8XI�y�6�^B�Y��x�Y\�p�5�
������컇�t_޿�q�_-��Њ
aA#x٢S�(ғ=��Mf'6�3��-���U�Y�+־���0p�7�w��0�ۓ*�}��ۗuv�G���6n���sL绳x���3 �Y��	��+�>kG@i�k��A�pa�2ئ��PS��O�%��;6�s@����H:|�*ň���i'f;A��^�������V$��������T�𓟪�$ ��*ɨ懐Z��Տ�H)!3�]�\q����
]�O��o=C]�4eo�z���7F�� �Gӑ[�8#�F�G͑М�yu>��#���&��j�x_�oƩS��=Ѥt�b\����$Ü�!����ðں���H���_y$s�E@P�>�`�p�$ ��G�4$�ҥ]/�o�9*�n��Y���/��(�`&(+�%���_��^�!Z�_�wDI�-��!P�h%�Ϻ�Fn�r&�z���X������Y�}~4�F	H�z�Ļ`�$R�\���Qd\A��C�>t�(2������y�^�=I6�Gִ�
\DL�z�C6��P�6 C~��G�S]�c`$�����3�ne�1�-� IMM�A�tρ���D
M�2�	:��l��
ea,,Q��ŉ�:=ԑ��fӷ��U���xQ���k�n-/��	4PK�����#{�\�o�(T�o?����������f���AlYzy����W�
薵@py"e>�Q��+�-ǁ��b�ew,�����=-xZ��ņ]�-���o0z��_I6�~����tX�j
|�o.FJ�C^����_���gB��?�������U�V���a;��`����R�'��-.�A�t�)Z��s��˗3�����A�l"��|
r%K��ԭ�C6]ʋ�&�nL�Bƒi��E���f3wH�C)�?w��bQ� ,Y�W���>X��7��M������jw=����?4WD�
��dxO��M���k�ˍ��M_V���������ysy������#F�#��PfcX��$j4R����a�O`'�<��������JgU�pz�/��@6 �nG�spǹ��[x�R��*@���ܷp{�*��WL���t%��)9�hBZc��0�Ai7�H<Bz�m�zy᧪S!�[��s�@Bis3nxee���񚯒MIR�Ȋ�էH���kM��@�Z�77�5�s������I`��4�D�+pi����uY������@�W;L[fw�������Y��ա�Aӝ�tѿ��`��6b�>��nD|Xk���k�ͤgI�8����� ���S/�oi�Z��v\�x,��K���@�7 E4��F�U:�CG\�PpOo�v�܄[�h��\~���>$�}S-C6��)�yf��3�q��C mႹ���uv:��7�W uo��~/a]��A�W��G����M��@E@̟�9�>į&�r�x�E�8�$1K�t���++�ՙR��ώ�*���]����N��_��i�F��2.��+)�0��k=���}58�Y�����*�Y�.m�Q�U��O�u}��o�l]gR�/(����$c�fB�&'�8��)Y�h,��)�����c;�!�9�����.	����+y��SSC=��5h��x�{4{�g��J'3����7�^��ɔ:1���ُ��*����>҈��M(����e����@qL\�)�@[�h�w�ܯ�+/�O������ؒ���5����p�����~��X���x��2�ߺL�
r��Aruc���X����K��ٙ<��ͣ����d�{���z�I"ef�A:z&�@Uyt$���ns`Z"����ۆ����3����ݍ�lv�ɕN�����,� d}�pC�������&��C�����N׻/.F�C�[�6Z��HS*��kF>��-�����������{M�gl����v�r�R�?55�{��b*���X"�]; ����1���p&:�o719�(����pm��:rȕ_�~2��ۯ�:__��ʴ甑O�ep����Q�#��$���h��U+ ������l�nWQq����H(ğ֚Z�^�j�5;S�f��7����?�+��:{䍺O66��߿�����+0��U��m�����}��s�`i@���X>�N�U�����ѡ�8�0���ƒ�����9��]�z�r��|I�͒�!���q�z���p63w	�`� �����9���Q�����F��:���<I3%tyrk�f�&��I?��<�
��_ؽ/����%}"�Z<�A�E�^��N#�h���ޘ��Ml���{�++/���OՅT�_Y�kH��(�(=dF<��Z�x�g������f�y�۸��M��WB���e-?��d`a��u���0�A�����$=��3j�_�_y���`�PŤ7����|C�k\w�����ǈ8p1��n�rW����C�CKbw�i�5D��V�|B�v%�ges����6{���[V����=��+��(7�pӅ�Kt�� �g؉ع�����#*-��U��c��k���|����[�d�[�IO��-�?��f'ʯ�����������J�3�#+����Ϡb��0��ǆ
��t�h1̮��'_�KP�Kh�/$W�]C�Y�O�'�+��$ӑtË���'NlLL�X�Zi��P�a b������G���>��7r6���]��u3��o,HWe��Sn�_]�2Vl%�@�~A�3��w�"3qv22�	���y/���ex}�֣L�hL��e��L $��Kc�u{�F���23U���@��)�K�鞪���P�G|xƃ�{}o:�v���)�X!W�6~��a�����l�R��_�L����3K&��ZkF�݁<�F��0(�K����������H��&�}#r�}Y�k�5��Չoa�0@�5.&�u����
w�
�OPs&&&����|Yn&X�;��
%��G#x�c��4�	�bz{{e�=�YJw����/A�Z����������F ��B�0I�˃���g_�"�y\�h��L��WB�X��b��K�DB��ȕ��7��~[-Xk����K�h�9�&�V�(٭6O8$�n\�ǿ��9��eR@䭧�L��������i�0��zǴ����D* ��K�I0e_}��	��ʁ�A�z&�����)��q�Yy,�J$~m�phO<�ĵ&�W��Uc����Հ����x=��{ʵ�>$b &���7V�#�l63-1%i*���� ޫ����n�@�T}�E�w�!C����zo�6�q�J�� ���S�8�`��7M����.؏��L�O$�/���3�]H¿l��F�No��A�Tƹ�����d�W|�/17Ͽ�Q�|=�����X�r�W0�`%%]s�V�S=�nQC���[�ã�[�k4V�u�6���w��	[GՋ���ä֚������Km����~�S�8t�453��H���������93����k��7�76�~��fZ������cn(�WW�Ժ��,B����ԷWݷ��������<�F���;#���q�pY[�f����g�N��������;���6��o-=�	$H��Bl��g||�r1A&���S`	�	��d׮�m�����.cs� �����&���+�^%��
Y�Ɖq�\�&��0Ծu�NglT=C���T�C�Z����S(@�g..?��ֿ<�����]�$ВL�¯���sQE��oZZZ����J�S��B8Eܵ���NM&�\Aw��I�w��yȖ��Ү���	���W�"�߬��L�H�����گ��r'�"���;V6;x�.A��J��倲I�z��!,ֆy�T��Zc�b���\�ߪ�R�+Ap���χ��S�����K�֘^��l�L�F		І��bP��n��>G�q�����{�æ���F��"w��g��o�]���#[�m��C��/|a>�a��+����\H�-�i�	�u�O����iHZ*�*� Ɨg�k��?�!�6g��"�"�����:e��'�����)rY�/��f�:�E��{������~������}����B:�S��y�~�+�,�2 ��2�Y��"��ӵ�ySl�|�-\z�����,I�V�0XV}x�')��˪p����,� o9@�y}jf������8&��u�+��ԧۗ�Ī/�mO��{*�u/�D��Z��2�G۞|��-�0��CF��!��%'?�u!#����+m��eg�65P�_U�F˗��������Q�Vc�P����5鑰6VII`b����XYY_��n��f2��ň��#�S)6�pe��,����EX��YA�f�2�0p5�'""�"P#���iN1��2�b6�e> �E��H�@"�	��)���d�K�/qw�>-�~��Ȟ�ma﨩u���^^p�}/��=�$�Ϙ/������5�b�60� ��l��ek?'_�fQ��G-��= 5��PuY�7V�?�m��͏ؒ`��EdM	�x����Dw�t� >�t�T{��$�E���;K,�>�-x���B�p=K{�����C{?0�8j�����6/q�����g�P�����H��?5ݗ8�)��~�2�,�=k#��q;�a���K�Pr��|Z������yf���7��c!�^��3�ךM����os;��zv�н�i#?���m?�A�'��������W�"P�j���%%�l2n�ۇ��u��;��@0J�k���$��E��op���@-�d�t�pk��~`�����/1<����^c���⠞��q@E+�Q���+�1Ar�����y7��O*��c6=�JB"�l��Y�S�@-H� ��!�[�P���w���z��(��Y�v������.��Si\�K�̅�8U�`bӌ�@��=v����yZ�~�ݰp��|}A/gk(###�v�蠲Յ��&��1~:*��LKr	�u�k�
*���`f\���y����\�͕b�X�ꃯ�bb��A���N΄c}�c7,U<H�2C�D},�u ��!���b�?���I֭�1��|n��*V
��a�k�]�Y�2�6q��A�/��@0J��
�������u�Fpr���`�K�T8�H��˘v� � m�q
���"!���5���8n��{ԯvY�?Rz��L�g�s�#J�Vo)>���r�]V�=�b���/<d{�YL�7I�W�7���Hā���A�b�����9n�žB 2�&H|���D��cC����)-�]�jJ��׺���X�W\�v�~ΰ�KȩyC2���6?��tK��V��%����M����1qq�����1��&z�o(�}Kd����/���ڣ*�:B���g�6��@`zu- ZP�H���k�\�z�<ގ�f�CN�z��Ý��ʕ��*��~#O��<^�9J���6`��c�N>}[�0�*��*����Ҹz~�o���o��YT��q�kiӶeVb/e>����@�v�� �u�1H��rD����[�3���h���߿PK�^�ZȌd�5󩱤5��V�f8&�=H�,!<�ɞ��;w3k���B��؆��`zh�;G�g�$�ذ�����D����I��������Nn�|�3i?������ʩ�R�Ɗ�:Y�|�{��K�s �@g�#{6i��{��f���[���^�������
���ȇS\������,@GQ1֤�K�������2���Hj�i���{S�/}2�h�YT����q�'��}�V@��g�ѯj5�5a��e"U�����%�D@mg!��%��^n�M{�D'�#	���Y���T�'կj��a����"sF�c:����"z����f�,%%���)�7�b��U2Cdbs���K��l���f�c��&�B�Ly�<9��F8Qz��m�oߊ2»~���>��I�6�*J�f�ky���p4Q,�h=q�!�r���&�(.��b\���yh ;"7�L��wZ�ڤ��5�E���٠��N��myu��q����[&�ZJ�Z�Wc�ZT ��cp�X�SӋ�l��pJ�Z�sVz:����o����}	Wց�QOI(*���UV��_�i-���n��x�nV��i�����ɤ�5322���:E]S�(�K��D[b��)���%xM��U0�do�lCX��|gdwOSm�O���U=�u�oy��]���/.�B���r�����ϵK�������F�du��Ӝ2�7�l�X�U�"��X�����o�������'���J�dK�ފ�YXG�-��ک�k&q���ԴO�p�bk��	�i�ڄ=�#�����������~V´H>��������69���x���ʠK��]��ec$6���wC?=��Ez9,���uvͬ�*��Q��NoJ�͌G�����
蒲o��U�q�O��f6��zH��3��H�.tr�ʅ�ޏ�Ԅ����٦���Q g�w�<�}fcc3��!��";i$�[��RNS�"���������yx�s<�a��1�0�rx��!��X����GvjcP,Hɰ����:�:�n�B�f��2���`��(�	Cn�
��.n ����[b��x7$B� ~��G��B]M�u��kȳ�\p�f��x����i�1f��D�:�u����oV�]�u����ݵ�{\�����y�J��>LUF����U:ؽ�u��2�ZZ9�����ks�����{M��Y�ҙ�_��)��r�	j7mC���4$��:��zOW[����7�܄C΍�"�8ȯ_o!�a�]ⶣ���!Y?�\t�۠A�"ԃ=ơ�>�+Q�>�+T�&��="��9W`�Y���*�6���nj��q�l�Ծt����-���/����&!w	I`L�A�E�iQ�6�o���x<����$!!����p��6JL��gK��3��H������B&Hk7.J������N+�PE��K��?~�0��ѭ�x\�=}҅������S����i3��]מ''�7��3����ӭ��ٳ��-�LC��X4]��GZ׮_��˓5��~��(&�f�!��tX�U�ș��[�!���<��>�f_�v �u�z�z���������lI�,z��KV��3�x֦�$���f��_����:e��	seW��&�,5����

No=ͦq]vD_�V�i���2#���A�Ѳ��M`	���7sҼI���֔�Q�$�g���K����ӍD{YYY���z��i�#>d��f=o���M�r���Q(&c�Kex3���h����|�5rs�g��o��_�]��f��ڮ���k�i�d'�Lq���Ϩ�o�,��p��۞���H�/]����5��3�3���h��p1{	8��	��v�V>>��:<�J{�y���a&�LЁ2�{e�����,>���|�{�<s)c���A��Hu���U���:�����tUYK�ߟ�U�E4�f�v+Og�t<C�Ҕ��Ѵ�!�~�Oo��Z`���x��<�}�2�����妊�ñ}�Y\f&ky`�BҴ��Q��dE����im-fdD��ib"�z�߾,���1%�&s�B�c�p��W\�1��#%G�c�R���B=Y��?���z �8�����Fi�)oiɣ�d�GR\���öp�����p�RǓ�p:���|�ȸ^F��n4�[�����.����T����^%���955�^�(@�1�ۻ�j�w�Nd���1ռ�9&�*K���4.q�/JIr�C+�ݴS?|�"�\����͆/Kq��{�q����.>4�
o\.�)�����]���~uӶJP�g�q�-�&i/�X��F�%A���=�ா����B�4� �6t&��䓞3�uP��u{)�3�>��so?���@C�O\i�s�Fd]Պ'�7��	S�B���B099ycվ���ߎoو�rT��>P:�TQQ��~uMW8exz���56&��n���3�[�φ�8����V���/:e�7	Q���;������́���㑴�3���y�,��@���Dih���i��+D�蘾3��yG��2]96��y��VB�6gQ�R0wu��G�Hb�b�N��w�Y��ل���Yz��o
�Iժd"^���oB��,��%�WיB��.j��� l�k^X���J�8#�O3�BMN�t\���Ƿ��}jf���8`������輟1��y���y;y�	�Xݐ���u��ϧρ�6�?��trQ4��a� � ��Y|������&	c�� GB�s����	�����*����%���۵!"$⭖�Ω��RÀ�[y��N�xT�=��[G�jL�iW5�CVϓ�㒯-�e�r������˹��ma��ӦBW75�������9�dl�o���!�>қ$����Ǉ�;S��<�"g�m��?뼔���H��Q������7����6����'���sk|�n�o����6E?�(?�:<��TK)	'n"q���(����;�↖��`����v&怹�ݸ����@��f�U�͛G��z�F���~F{��O�RUo4^Z[^�e��!���|:/q��1�v�}ė�
��,`�H�_#��h�I�aU�����P<&�����I:M�o��_x�����By� x�Bd�&R.�?$K��9h��v�����Q<M�kg�\r�.�g_�m*��V�_���+b��p�b�bP?��{��N���Nն��&?��շd���X(,J����i�!,���X�[�8.]6�?#5��.?��@V� b���+0���&&&�ݯ�}肍��Ӆ�/L'/�,����j�{k���-�h������|
�?�����s����������98�Y��q��E{g�F��2{\�wD��ޖ�a�L}w<�����(!�ޛBR���;�W���3R!�؇�ñ�&��X!�����w�}�?�(��u^�9����`�3*2�@��S��6}��U�1SR�#?^\W��8ꖨ���~��yk8�����K�~nk����J$�*+�ӧH$�",q��v`af��ϟ?��E����6l�*B~Z�_Ý(�dez%p����*�ȇ	�k�C����1E�Ά7Ȥ�@���y�����_�����GN�7y�<��IQ��z���_���w�/�OZԎ�$U��(�%%#���K~��E��Dh�������ʦp*�b�c�t�W%J\F�y6��pO����Z�ڔ��J ����_�����)�� ��]vwt��ƥ6蠒_+Rp'���Gt��)���/c6H�N�a��`6��W

���3��[=߿��x������_���d���]��a�|1�G�ٓwg�q���C���"�z@�xMeE2�&x��K�(�`z�x��P��kt�5�l&~==�N���ź�����gƾZ�y�J~ڢ�g���h�
c�9S��W�6�8�7&A��g����<�?R��'cUWf�w�S����U�YxyѢ<6F�?� �G/�}�����R9�}��Ѳ����(@��]�Й"��TI̍��7�P��0}V�T�~8��C�����a����d~�]���YY���y��y���`}�����M�|��gcQJV-��='�yP�����j��;Z��>�a����	R�[�;4Y���%/M~�����dKxf�����wcD��`���E)��^��-�C.��S�ȷ����<E@):-�����V
G\U-�;�'�=��Z��D!,����QN	iizI�����S,��?,�mZs^�(���aS)*���~��i���?��3.�E\碟�u����
����0MV��+�؅�SU�f���?��6��V�{�RO�4��A���]7��L����������8;kiV�p�,;A�-�F�rp���!6��oibS��1�23�����ʓ�bF9^����Vn���ƍ9/Jf;XI�@QQq�/ �Po3>*�0��`�=n�777�ߣ٭H{�{JڔW�r�aװ1J�J]�6��1GG�I�Fru�J���1�S��c!��� =I�Wr*�x����SNhr�.���7l�^<jpY�9ށ�ևþ�I{?�^��Z�=���^o�0V�?��1���ݭ89��o�x��_;��rQ��ݵ�V3A<��x֌*aƆE=��7X���{���0OqG������g���+�?U��U����Z�z\^.s�݋T�x�\`
�[�#��J/��C�d�>���޻܀,�������C��-�����.5I��,����5����5���W���r��.ЋC�w�>��Sq�ϡ�-�;Z����z��>'<	ʖ����ߔh��&���̿B_C��.�.�v�žt=L����(0UU�U|ޫ��c�b���ﶗ��P~�ɲ).��mCG憄�4f���QNVۣs���Ɗ�nn��3�P��Y;�Y?!����9��J�&�0e[��}�C%�Fô�+� ��,.�OD&���@�nh����x�~(���m��4��'�(����s�h�%���z��3ظ�_�a��/�P����2gIn7���L�8�L�;R�`W1D8��Ow^�B�^ܥ{�������m��9�r7���]F�^�k[�������kRѩ'>���}t?=ݵ����������#rӖ��҄����˴U�#Q�Yg��ir��
B��5nLT�ޝ:�3��{C^�BAA���H�~�75��^���f'�Q_O���82�Tcp�ѣG���nS�R��5��c+�GY�����_���
�4��u�iK�i�5>�./���',��η��g<�y��x��#[�F03Li�Ԛ�q�i��SCv�#�IP�vx©���H�X>K�V���������~��H�fw�6��B�"nߩR-�]4"�u�s�&W>�!�z濶���%x��N��p�O㧑b$���$�Nuv�I����˅֗�/}zF�?�֍���#ٜ��q�k��u��]8�2�612�9=y%�R�EM�U�KM����#9 X�U��n����������D���FI�ذ����O���͍zO@A0��!E���JA\�W�5 8(X}�����v�V�Z�`�����l��Y��}cܭ�K����S5��HOƛ7��^3&l�Չ#�z<C��v"X	<�F���ng�{M�מr �����,��{��r����e�SL����C���8��)K�Ɋ[��N�h���q�r�U��������NʇG#U���O6����%�=����g ���g��2f���b:]���:e�,��˹�m�
k/�"b�D+�$�QL�������Ш2�_A4}g#d�0�=��uo�ex�����(9�A �c��c\Kۭ�����zᗝ��ve�%vޮM��ݬ���Iy�w#�����1aA��:!�3�Mu����#^mv�WV�jR�=�ْby�y�����JzŰ`����i�:l�'��
{ӓ��u�M�R(����׻�ύ�2b��g���,�3�`�m����p�7;�!�.5G�ns>m�H��1s�߳�J��&~C����{���3}�1Guаz)!T!
τ�gr������!��1���܀��@1�B����&)	����ܲ��~���=jN�YFo���c�V]��-�y�f*�.Ѹc�F�q�Q�S�G�I�����elj�=�}q�!IS�ݤ2@Y��M~	_��&]kn�mg1�O���$����d~��2�ޜ���J�Zi�js_-~4TZ�U�-?1]�{���{L���ü�a#��f\����;��o�*���CQ�F�8��:a��E Y�gAK���J���4�����Pw�z�NM�/��q�%\gD�^�I���=����\�_�`�n,�&�*>�HpΓc�ݰ!?2�{�����~�ߡǄ����	�#�v��/桉qwr�}S�>��J�G�cb��V���qT�P���|�`��"�%C�2{�d~c���'O�p>���\嫴�UE�����QI(�M�?�n�ɢ'���WV0O���S�c9	7�%���=��/n��̒��b�;��qrw/��Ö�3x�N�ñ8@�F�?H����T��F[�n�FW_w�v�]:${���Ku���'��8�dc�+��5�9h�w���e5BeUF>[�zS�������Um�0��/��n)6D��>��k�M��݅����r@���ʕ ��\ȠNj,q�Hś&���NU���W��RP�hǶ�{��6ez}�?��gC1���X��	���:~���"reI�K��(⒒��X�řъCZ����&�\Y8:^���9�8O�K���Ki�##�^�7��1��۰�Za�p��`9f�%dx�_�9��%��BP�@-��fZ�7��::ư���[H��>��gz�70z�Uk�:k;ɨ��۝�>�˿�u���1�fD3[�v8�ǋ�}����6�=M�|T
(���/���(M���E?p�{C��azQ����I��iM7+�i�c��/S�������~�:"��=ӋXl>RA��K+O�b-]�� �j�l�=Zl����b��n(`�	�1��t��ߧ蔘�����ﺯ�<I����-���U:�I�]KX+��ǿ�6��PA'���r�Ҡ1�a�����Y�O|v};-\~8�!c�1�,�U<�5�
۷	H3V�D��+����!!�&3`���ww��7ǭ)�%�zeN}���{���9�(��� �	��O.]-�9䖔�z���gg����/�QH��a]ӑH��a{�:�Oָjz�/ZS��5���D/ϣ��ͣ��"�p��PI�G�5��[����8�*x=�%f�:�Ъ�_sT n�!�Js��e�O��Ki�IJ&V�<��w4��m����^���7��N��"�d�m�����V___�2�塈V�$D"zK�xN��ꎳRk-[z��y�ԟ�ȁ1�=4�K|$�����.웳������W<�Ս�	���i�^��ؚNδ�aEV�ơ��6��u�#�\���T�d�S����BBB�#�x�S7����Z�Ѽ�f͞ �$7B�.���Y0k�a�������bm��rB����@�.4��h�=�/�?��k,�V;H@���U�����
�7�N���ro%��%oX��Ic"7�_��%�}s_
wLY_n'�ޘ���w�*����"��|��*lw6�����K2�s��$V�^g���{z�#��UtvN��a�����JN�I���'�<��rf���.Q{{��
��&<�W9��9kl�]K��@�|�MM����h,��Z����*�:!-��T:�]�^�����S:[u����%Pe��b_}-,Z*yV]!lnX�|�aC¸C��N3���u��89>�c�G��D�4A�Ͻ���YV�GSk�D�2Wq�3�֥���W�/�QGH8Ͻ)ؙ̧ۢ�A9�#��j��+�s��::�p33G�i��G4�S�,��|��qMбw�V��=ƍ������}�FshfGo�x�8ϣh����ll���
�k1+�8$���Q�w��B���!��� �D�H��y�}i�����������g�bn��I��dHg�G_���XEE��s]%8��C����*�:�ЦJ����K76�o�ݗ��qt|v0��E;rK��As�������X�õ�4�tpQ�\��H�2 _�8���ks�gr0���u��˛:���O�}� �Ǉ�h;�_��*&�|/r�?x��J��f�[�H�-�����]��J�s�9-ͪ��x�~aq�+�U�j*�ң�,H��Y�o�H��|��d�R /K��C��53��x�P�y�h�Ac\i��� 2GԹGp����G�ʺ��-�O8 ��h5�FFF"k%)��:& ��=�m�4�z��ٵ/���K�����w	8??*y�5g�d�6�@!�?ܒ`��a�¢������{k�r)B#|m���T��G>`���������X3��'~�͂�o½���I���lg��2h%��g�9J.zm%'�ĉ�.��A8G��ڿ,~��Ȋ�iMի�{̕s�^^��(�e]b���l؊�-l�M���q�ϟ?��<�Uxg�Bpǋe >�gr��O���cn�ݬ�Y���_����+~��<6ovg���}���y�`g�j�D�j2�Q�x�NN]�y��uZ,NAu���x��\ʎ7y��$(���L4.n���邺+̵l\��)���&��.b�D��p��W/,�I�
B�}b�e�˯��87�!7r>?7�K7i��dC>���鎙aE��_����q�!�]�a�֌��J��̜�_R
�k���]Jqn^e�q�ew�k�;��9��]�5�3p��a�%��ݐ�:^�s��꧖0���e�g�4:�afJ��.��^�0\k^�H�l�h3�H7�����y6h�y��6�m�6�����i��r�VGK褉bY��7�ꧣ�|��u.Bp?��	�~�m���<F���;L*!�$h�Wa�.BLXz<PS�)���|-o�R��OM�U����l�[	�<`c�J�}�~%=:�I���			�#�:#!�>ZP���Uڨ^���Y��=�#:d�9�~|��5�d��M�et�N/�|���spp���?T���bJ̼9�.Ƈ@�'������T%C����Iߏ��xg��7����Q)7X>_^����}��mKqv�߫]�e�+���-�m�ܪ�u��	|쩒�ߠ;=2�#�ڀUڇaT���at-S�IQ/&k]k���t���5�~߱)�OS?��������v���4c/B{�͝<'��ͷ��͙�q����Y��,�@��7��+��iZ�A�$m�����$��}.��(����4���ƎWYEE�o�@�A(��#%b�hl����\�����h?z�P����ߝab���B�br����G�h:yrN���"��r>��
L��s)�%3�]2�l�#q��[��7��u�C@
-a+2{�7�oF��F�T7[�(�J�*���^�D��&��w�[���98����F:7��'e�p�ʱ�Ҫ/�N|��&ʄ��$�Je�9�a%����|W~��%C4��j���Ŏ��,��}p�
��I�7�n���˜�G@�y��l� ��<��ߚ;����
昲M�^ڡϯWX�ήP�����e1m!�Bl¶?>����_ΰw����[M��5��#�qy�븷r\bY�t(�E6��}��Kh��tb�Cܼ�l�T�Q�S�l=E]ϽK�#Cv@�غ�վ�-ed�-wPy�)�\3{�l�C����	��������~ۚ��AGl����,�B�_oh�i�Mr�&+:���=9s++q��p_ޕ�>v��~rZv�&��Wܲ��'&&�k:z�5�[�f��v�������k\�9pYݑ)3�b.	Z2z�H�ol?
�8��M�9&�d�R-/E"�/�,�;1eB}���b����7����$�2֧ty�����^dY�Yo�_:�W5��XA�:*�|����T�M�V���i�%�1��H��&�AP_������ijxA��wG\�?0lns%>�N�H�G���^��X��چѓ|�T�H>�x�}�(��4߷�tX���F:U��=���X;���J"���?���qЉw���p�[<��o~!�n���+C~��t��ҟ�� =o���U騕�ö6�v=cc�5� U���ls"l��h��"1LK�)$�`��g���lGw��v0W��g�xP�4l�B�l�Z6��1�5���`��u���l�����|�yT�p�|&hZ�K����}���,�7�����m��$��A�<*o�8��P�N���L���y�_N�W�.�	pq�w�[ɾ��ҽ��u.��������ۯ�ڑ�V�����fsK7����و�s���+�[���5��|w+�Ȯ��0j5@�Mf��)����9�Q�<&M�D?>�-�'���{@Rb�	\s�ɺ0�ģC�c���	�R�A�o!.*د||�a��k&�F�������]�� %L�E ��˅��;�{q:�/~{�������Q\G �>�|��v�=9y�[�2c4mH!g^"�Z��y��q{?�1����R���}���o饒�0S ����?�97�g|j��0 �)6�PY���A0x�J��1�P��{=3s�^��Q�s�[b|�����7ox&ȼE.
Ժ�tB)"���m,rѯ])t�!	Pk;���o*��8���CCl<��"�r���,�tb�%�����ښ�QYU6�+�\��f��\J�pAh B�m�Ep�+3Ff���ww8���U6�@Q�x�&EF�)�+E���ս����b�o#Y��:�E �F!Gz���[��3��{����'U����;�Ahww���>o:F � r�5�A�JFK��X"h�6����Kl2-� �˛R�{w��T���ܦ4��pO�1k�SZ�y@[��
�6C���@�|�څ��ì
�����߫9�/P���/�GF�C���EFs1ՙ�����e�nvuuM�����9�#mc�����4�|	0�$��W��~�p�t+�;���.�cq �uʒ��r���6�^h**�hBSL�'g��ɦ�_*������4oTx6Z�Լ�~t�Ձ��1b���d�W�s'�ܪW�)r�렚̱4|(��m I0���zҠp
�oB����d�a0q�����}1�ۋ�����=	�,�S�Ճ���G�c��"h����M'���?k]{��E�T�۹>�Q�Or~�薔�e������� 7��"7��bȂ'���f@��k�e��p���DT�c��y����鮾���Uz��=\ ۄgqT�W"g��".֏�B2!L�@/e�)(R�n2�B��y�j���������,禧U>f�mx�ż�G����?7]e@�)�ߏ�"��r�'ռ�p�b���H:u09�'�Q�/�ң�m斘����+Ę�:'�~����k\���"G8)x7δ��k��r2R�*ҡ��2�?K[��byӯ0T2����pαC��<�&���H]EX�� ��Q j��N�ڨ���T���Ϸ7�ﵵ�Z+uP�`"��-�����M��t��U8<��c���ښ�w��1	�#2��u������?�F���!$@k�Oy�#��v�c�h�ƍ�����fR��Aǎ�}	���SvG����V?�X>L�,�����<Ah?ޖj6`�7�8[9��ǯ�%`|�vƀ��{�`$^5�����H��p*"�j����M��9����b�Ҵ������q۴%_9���P���*�"� �;^ai`l��xx:<��KK�LD<�h��%ݽ�˖DA9�en�G�@^R�F�T�ik�>���;�O�eX8ER0�fM��JR�k@9qD���1{Æ���2�5���?��yu��p���zW]X�x 3l#Z����#�[N�����`S	�;=
��H�#�dqVI�e��09G�,�/�r���k��Ɲ��ό�9�Zێ񘔣�u<���g.�J<4ֵ4kJM��a����6��V�trN�HJ�?}�pp�|?���E_�T�H�'��F� =^_���LMM��z�����K�6W0�����iK��/�
�)dF?_q@�|�*27k���E{��5*z���c!5*�e�͜hR�Q��,[{��ϸ���I�#:�<�)�0�I�����d���?C;(!}�H�SzZ�t)��w�����n&�=>���n�G��b�,����Mh�`h�O���x�"�[Y&t��[�����U���WJj�
���؀	a�(e�Y"H�`��)͉����iM�W�G�Q��ʓ�_#� Q�{DnsQ s��ډ�''%e���Y�qRL{��U?��L��E18YY�d�.����Q���Ãs0gՈ{�S�ޙ~<��~��O&V��w�Oz%???���P����h�Jr��O��� Gb`�"FJ"��8��0�9���U$Z'xh������W���<��Khk[��G;�J��I�Y��׀s]�s��~�֝�{�щ׏+�a�LJ�Vz'���u-�*{�6��a R�lڅ��ׁЏ��m��sp�����IM'�o)z�(!�����rS_�/�/�Zk@uoJ�uo��l���F��	\���lw^X��(Y���	���i�m����Yt�@��ˏ�1E�MU7����ͧ���i�=ĂIS��n[���iσ�F��Zzd՛&m��Uo@��n7���6��q���h-����������$%��e������(���o�#{�a�LT����%$��3ٗ���uE�q+����y�����[6� �5�S6-?�#��N�N�FFF��rH�:�tb}�qꖽ��2��ξN���$̮��y��F2N^�\L�2҄֫����S�Eykˀ�q�{�7vW��u��6���G7�yyuk��M�҉w��痋�>i�;��"0���pң@��4�ouu�����oS��m�ngg�},L���k0ZI19�/]7�E>�}h��h@��ÀHn��x���8���;�Z��[�7��拾�A�p
G��x9��7@�m)�O��aV�ƭԍ���\Gɦ�22�f�M�AL_ƢP�y	P�&���@�I]Z��@��1�O��mti��]�V_7����� �7��b�q�C�M1�[�5��.�(&=p�0)aȕx_H\��(u[ ����0�MO����49�I/�[Z�줻���Wۉޮ�?����o���3�6�^�|F@��%Ի�������Ζ����	�sg�1�pr~�F� ����箮�Q�>��h~�:�z�^��
�m�DX)7#�,�/��;^e?Z���p�C��,��g�G��'�ɇ��o�fӮ����[U���Y7�@:"�J%��[��y�4�JV�ݣ���a�I�M�������(z��Ǐonv��\���ꍰ�m�4��u�ro��~n��s>��lTxlL���iQ��5����R;�V��녺��Uܬwl��8"LtҖnz��~�3��P�2�nL|מ��F�X92��|�`c�5�����y�/�0��wKG�fB;d�;`dݠ�����0l[�D�9�Q�NЭX���b�oT��^RR�B�ɠ?W���{��?��;�F%��^|��x����J��a��-�Q
����ȋ��-�)��oc^~���zo�Kt����%r?[�J��A��:���k�!�[�G��]N���,C�ӵ��&�O��.M�N�L�Ǚ���y�!�������z�*	���~n+�]��_J�~�wX�߰��\�0�L��kp��Β��q�b��MX�c[�?�l��环�髴44L�C�-�@-������
@B����W�����ă��{9���}@�T�L�_��fh��芿hV�M}Eٱ%����D������O?s^$�9l����J?�4�N����o��KBL{��k���*?#��\���~���R|L�^����{�?g����ׯ_1?zz+;$��#Yq/�^���߿���j�T�+�ܷ0�o��_s��^�$"4�@����|N3���y�^������q�r�9~F19�>���N�ؾ@ګ-S7�]=�Zd���R<��= ��$�JI�����R����b��"���L2N8�~�lJ9�.V��a񉮶8TO�SG�%����8/1B�t���1����jU�7�bV/��q�r��پ�kZ����аR����u���80b�&?~��~Ex����Cd�r4�Q8�zZ���h��N�k�%n�R=��q<�/S��$�~af��`x%7�����&�0�|�2�&z�@��=�h,f���B�N>�����F��f1xؓ���c��MX5L��~��a�쵖�r��>�uP�|�p��đ��?�F���&M���Ԁ�ո�'I�_���8
}�T�Y�}}Md^��>�\C����Ι��ݗ�(,��=ϫ�~�"*߉<xr����c}��5�������1�~��6�1M�����s;�!��o~!�wBv��8���4N�Ԇ%��=@�uP�[��Q5���N9%N����9��\X\�����1�Y�V�'���t���F�OBz�gP��k�AE��E�$�?�K6&d�+�._2�Ӎa�c'�8���։��R��?�}�h�i?�v�3��跳�=�w���3+��=�	�؋iKW&E�Z��8�3��)���4oW�h��:���zg�k�e� )Rw�t�;����AZ�L셇ICl�ư��n�e�d��2�P~�je+7M���w��Ҁ�?�XE���
��fV�Υ�?� u���8�4A��g{�S���!r��V��)����
���j�]��c��\����ALJ_(�q�B"�<���8I�S�D��	sQ���[�^]��=�2Ģ,����I8��C!�n%��i��xt�qQ�ǡ��dU�)G�hR�{6pGPC#���O��\�?H�"���eH$�~&�)�i>3����'*�˂�����ᆝ�vz�a��/��^@Yl�����_}�GX��D���#�л���>��k�O���r��-�A�h$2�[��8������Xeg�9�yۨɇL�?�S�ޒ0�Α-���:_�,�> �s�CbE�fb�CP���[�,���3�.�I��T&���:��Y�0���j�Fc#��QwA�pC�BK����%�����+g�&��L�P���O���G�۰�Oe֐���h�WUQ���J��ҹ����I���v8����RRRƨ;N"M�_]�d �1W����l����
)���$�)��bDF�dT�c��M�G�HnR�
M�)���K��YW���V����}	1��mQt��2o�.NwYz�6K�E�0�]��׌����\���āz�TH{ﮍM/�,��b���F����PN]=��)���
;�4
�f�B�Ȏ�g���"��&�k�􄓮��yޘ�3ov3S0C�.�Z��Xu:yte<
1�}^n-�ʸG�d��T�a�Rm����'�ƾ�>JY���A��:�]�Ã��ģ�<#�U��fߙd`��D��߁�:������j33�_i�S���b��R� ���v�nܦ	ӕ���Ȱ��׿AuJ���O���C��5�t�g� �S��a������A+����n����Z0���1���q�a��ͯ_�m�¯m_h!jZy���h��>�v�Z���{S ���H������{���������h+�A"]j�����5����A����D_�Q�&WX�#|�y���e�)�?=9V`xxs�V�{%�YTL�9A�J�j�T���Щt���&�gU`0�6"ufK��y�-z�a�����W3����,,TŇ������h�ʐ4�9��E�)��,�T�$�A����(̈́Uf����&Ok0�܄ʼD������0\�ၡppF%�mn�����%ɉ���X�B־;N}���Ӊ�S<]������d��ZV2<L��NmI�@����^�'����Dܺ��u�	�)L8�'׭0$�@�^���}h�yTA�bA�5�c�U[
;qa��>3������:����Jz����ſ�f�%</e��ޭ�[�-N?9�t���7��FWN�v7L�%|������p��kɨ~�gϩkx!"��H���$V�ۅ��8��ʊ����4ܔ (��)�:��!n*M�	<*L}����l�,�Q&mb߽{�%!@��;�����,1���iv�l⿰HFݢ������
)����T�A�7Y7�ipΰ�.����!C�D1�Гk=v$k#�@z:@����s��E���PSni��*�I�d�"�_b����NH k�~p�����0J��:`0N�C�T
�����o�T<���/õ����É*�^_����aP�I$9��X�_ːUL�7���2 Rjjj���ޤ�$pe*�h��P#9����l�xk�>�FP��c�@�X�������)E�֎P� &�����<#+�ɕ�,�#�K�P'�c��a�_��������0�Bѽ~}}}ɪg�Z��V1o�7[[�b�%0�I�?�xhn��&������Im�`5@��P)spkO�	���?W�n.t�����hkLҷ��Jh޼�O���l�!��5/�6`��"d�\�Ŋ�"Ѯ@e��I�*��0W[�4!9���7d8��g]�Z� �2j�K�܂B"l%2T��A �o�y�
��W���j�P�V��MĎ<��"�p!��{��wT��p�C��Li=z�ͯ�ŕX4cQᦎ��L}��	pW4��*aCP�|��\�R!�Y?�����,Es��Ǟ�BO�Q7Pa��R�^�Oc+++�ѯ�b���g|��FZ�c3@�Mi��� ����z����&)���b�	��K��T������R�j�"~"���罃��������o�ңa.�XڻK�e.5�Eύ�B4H�����W�Y�1m'G��Ɉ�(+����]	�������A�鋸�Wd��}�l�N�|h�t�L���������;n؏�C�����J��Q
�*jj����v�!G��n�@L�����D����o�;���l�w�����������$矇8*vO_��g�M�7ȕ�s{h���B�*�Q,m`��s:��	$�͑�u���?��I��K�	&�����������N�P�@��P�Hl����ױ����6��5�k0P�/w���h��F��L"}���KB� "Yi��j�<��eAn��d?�A���d���	Pnؠ#֬��od=�1�B�����4��հ�Ka��a���	��ޛ&}���>�y�B�3i3H�Zh	n�M��o��%�ݿ{�h��RC[{���(u���cS�_���[�6�fՌ���;�6�Ҳ���,@��!�LiP�F��=�g �eR��6U]V�"*	�'uDU7�"7����"����Q;��q4��eF�����$�%H����Vҙ�"�l�Cf������Q ^+y�iw�>&;[ZZ���8�#YY��4��h.7����$�K�
��o���:zv�c�������v��%@�R��D*�Hc')��jkm��\V��d�iDu��p�jz�6 UA�S�L�	�d�������@#U��U Dz`�jA�34��J��KO߃8}�Œ��u��,:=1C6�@J�����S��	�y����ۇ_gf���zsN��y�['������ȉA���y��V�˴JPmm�KA>�,F��}���u�7�2ϣ�7��e��g ˌ�UIr����ך4�6��ԁ�Ӳ�M=*KoÇ0�	��`�8o����93���f�Px��P@�fᰊ����az�t�p����NpmW3�y�^%O,��I��cvcU��5�����d�J��]b^�[� z�Q1ۻS�;LZԘ��=�~���F�6^`�U�o�h���Ei��p�V�u�����x�!	�|�!��f��3O*��?��WT$�-�/"%������T#���)���X:T����c�+�ʣ᫪�Y�ձU� ���
)*	
W!�ydcgvVS�dEh�����c#	n-�M��9���.U�O�^ ^��e;�N�ڂ�ː6�� ү���V���!vs�r�aTGx�+c�=���ʬC���ݻw)�~ P7S�
ȗg��'w��
�|�#Ľ����m�� k�WىP� `Fԁ^�zk3���BJ�?�"�L�4�׎�Z��F�񭐿YSB;7߽=��@ZB��*�ъӲv7��ұa���� k��GW��5p���C�L����us��|`��k��j6p��Y�Q�����eƦud�ǔ�a � �J���{^�"����rk��K��<�:����r7���E���2;�X'���B���gV��w��7F݄�2@ �e�c'N�5Yg���f<�(��]�?���{؊�0 s"�f�K&�．DҞ��q/��$�_)���!A	Җ�Ux���]��3�-,,��C��˻RO��&9TaE�"̽eB=~��>����wi�?�&8������6����D�l3J�87Pz�4r���R����J�\l��?�&�| <*s�5���
|�G���p$7|!#�!|��˗k(�B�tگ���
ܽ�V��5���юX#�o���t&�Ҭx�}�6��"�P�D��>u�o`�%�P�xڡ"3��i��t�ߗ�ߛTd`�1G�2���
��/N�1�wi�=@��2��[��vgy\oD�j7+�-r���O���{c��̰�(w^�nB���"����z���wҖ:��|��
EYLǶwR�m{�/sd���=��S��ӧ`��0(�u=K/�k}��9�i��Ä���,�k�Q��.3�X�<�F�b��5��Bh��3h* /aҪ;��{�X����*�� �q�N�� i
0}Ǭ�{P�p�׊���k�^s$w��5��BC;ZZ�,��^��ajv�T����@��T��mwm��6��
@��U�(DK`OO����ӟ�0p�	��M�\�>l���+�s[�/��8���)��x����������
��b��R�k
d�K�%��C@X�����wwUH@���W*M5�s5�vs����kD5i��M�aQ�᭙ ��3�d2<���n|�B��\!�肿�[��z��ˮ����-Zy�����K�wp��������=���������)� U0�/�/ y�|�`:;n�nX���qU ��<hO~��9W��o��M��%���o���X=�@��������w��EU㹵�����l�(�]�G���sp��h�aK��*m�yܗ�H����"Y��-M��y%�\A��J�
{ޙ�Gw~�TT\����㡤�Lٯy��:rϵ���nacå!�����*���/�[!R=(ӕ@γ�	�c�Td�0\�uo��&*)�}@vh�����8��� ���J%4i��Ѣ#&Ϡ���ⱶ���Ťk,��b�\T��\Uݯ"��RzguoIy����Ѫz�Nv�9�(��V��.��v��-���.)(�?�%�W&1�9l���ێ�tYUQU�����n��4Z,.�ĕ}�<񎞟�~�Aqb/	���@ݵ�����'��!��K7d 2S�x������3a��g-d�%n몍�����=h"��u �6
��Io��ә�>���gk����@,ŧiFs�Q�]�38c� �Sh9f0�xtU!hߙj�.}�1�bP����l���j@����3�ۋ}Ċ�F5⎞�Q�$�n��=E����vKc���N���Y�S���@��೘.%U��*��
'�w`pVtb}�c}Bg_��,1ȁ^jw����r�1�5l��ָ�����	�PT*j�������/$PN���)e��3Z�=�O��Y���5<�^l�ȧ����?΅��0�gψr!�����7._�����Q7O���K��L��g*�}z�}vS�̓7J4��oM���QS��P7�HSS�!s�E8�{�1�K����_I��%�LE��!�j~���JJ����6H��j���dX������94��M�'�z�sN"��=7h��Ӟc�j��*��? 4]^^V�Z�����������������a�w:9$ ��H���ď8�S�`t�Ϡ�AݫR���&� ��z�$(c%������?����bׯ�u! �
�zƻ>Uѐ�o���� ;��4io��u���rm��L����۾� ������������0���L�%����xp�zV��Wl�����lm1�Z���'�:	���Gr�\��&�@9��Ĺ"�����
'���O�y
�pT_+mG^����~��3�d���J�z�$W"t�,������Q�ͼ�_S|8��sp���VIÁ�.�FpW�I1�΍7�{���z���F���P��m��TUU[�Zִs'xj�Ҽ،|�{��2P� s�����p&�1+�_+5?G:��߿W�;�>N��u��k�N��뭅�8�M��a�n�W��g;�]�_]�/+-%Gm ���i�1�sNZ� �?�9���$^"n�»*���̇@��F�F���H��Ƹ63]j�df%�y�'M`HW����B�7a|'�!�#�fl)��uw}��E�ϠʲהPSԈ�u��G�#��M_cjjj��_.�i>��Yd�*�����@�Q��I�� q+eB�j\�K�4M������o�g*��X�8y_�.|���0#v��g�KgF3��)�0��d����:lH���b��$!��i����z%�����+�ߝx�l�v�l����������ޒ�hx	����fy�<��+9~ ܜo9ݨ~o+Fda	gv��w3��.,�iװa%������{�p���xZ�)���HBY�,-��!�!K���(�=!�p!iȖ})�d;c��������}��z�{�����\g�8�j�|��~���k�?��0��3ݞ���:M�c1�ͪ�W�5U�`s�\'���Ó��� �L���N`V�Q��x�׿�93|'��,9��n�*@+���	���A��#��拞��FY�y����UȺ$%�Nf���>_{:�A���ؒ[�LBD�p�Z���ԝ�ԗސi�E�ۨm�)(�*qJb����IY'96�Ho��I���*�%U��U�WN�x�ϊ�~����L�^����[���,a?7������׆���}	%��9U��̬)�I+]��gzz:� ?C��+���vI[�A�_3��uzG��e����؟Ir!߃�/?����)K����e\sI�7�77]--��g��5s��pQ/?͆�՗���m�����>$�thg�˃���x��h��ǩ��������o�(/���m�m{���;Ix��֫]��!����?o����F.Kp骈5�[�cx/\�6#�^`���񫛟>���R���O�v,�
d	7+�=�Ƨ_�XL��P�Y��v�����	ξ�Q�=��͉B�q���מ��ݲa^	2j�ǉbT��f�tP����5S{���e�y�@���Q�]��}̸�{_]��y���n���'����|����'w<��c{u�yx�iYD_���***FS�0E�����ֻ�+ٌ��8I��ғ<��}�c><�7_"��%3d&=��t�"Ҏ�Z:lǒ���ʤ���%x�|�Bt�gwh=�h��v�i�Sj�n �E��]]U����I��f��>9�<OL�V���o=8� �]׺��>������Y������F�����J**�E�%YY�&''?�_�v��Bbu��=��¿�<���/_�������4�T�ͭBۛ���-Ky-w������u�M�eq���KmD=�>:��:�O�|f{Mi{ˎ8	L���wz|�|�1�h�$o
�N����k<ZW�8�����x�k���tͤ��"��x�O$%��)��/�\?T����<�ȝ@6H�̗�~���h��i�g�K��r
W�'� 
�Q�� uhl��@��w}mޣ�J:~�����~����$��%>j�䉎����y�P! [������K�OҮ[�tq't��z�������=d���}�0>����fj����A��B�z#a�ħ��3T�8�������M���%	$��yo��M�Ŭ��
��>�ΰ���{�(��i,��~bD �J�Vɢ/\�1�{7�S(E�f��q��H��M��W��Ǔ�EX�$��p5x�-�/�(�ο�hO�N"��|Q�/�.3в��Y-��ć��i�x6wS�j�.�7	���~¿���:�$�@�'DLd���q���x����V�����kegOz?�]�5����Pk�$O綳��b�[�N_�}�,��%(S�4�����I�������Uފ�92_�l3Ց_T����u����OO"�L#�b/j�512�z��0�iN'8�2�dO�tR�ߨu��N`���;^ �4+#E8��ą--9�ܽ۝E�hK�_kQ"E��#��Ρ������KR�V��d�g��� ���޿�cs}�ky��/v�b*bL�W�׎�����ʸ9:YwnS�*/z"�~5��u���^��Z�բ\`����-������<K�oPZߌ�jN�ˋ��R&����UPo9�ӽD���G�s-�$��_;�C�����E�p��2eh����`�We��x���L���h�5��pV��e�CI��d���'_�.*�Y�Ծ_������I롣�܋��/$��kdX,J�=�5��/boE�г�"�<�ku�Rb4�׬O���O�ꘋٔ�̵oB<���d�vp�3ag��}r�g�H�:::��U�� �y�+�b�3z�?BO�ٷ6 ���������ϯ�z�'Z�u�mc|�ܕ�N��xX�fq0��Ys|Ul���������rs�r���{(�)��\_h�ِ(�8�K��$��cy �&�-�cN\��ٳ�s���z�	גw�Ђ�*|a[�J͝�<]�.2�����|�un��c���v��U���^���z���w��+��$_�������l#��޹s�Ϳ�(�G]]c�2u�g�ڣ,<��BG�u���寖��*�/�a�a�puO�z���.f��Ƒ�m�'�ђ3�#&P�/���G�-[��B{���O`��!�/�=r	�
`)^��xf�/@+aX0`�.�z1º�Ƥ����f�lIX���GF`->���a�OB?9��� i
۽�~d�}s�`���<nɘc���g}&��@��(��b��O�����ώ|�౔n8���\����m�.,<�h�z�)C�=�:�<��E���D�|��مcm�Ш@92��A)�&�R?��ֺ�|"TJc��`V�⾄��6mÈ@&���Q�����-���ڔ(� D����-����G(�ǓJj\��Ɯ��٬Ah�"�?����.Nz]����W��'�����$��gP���>��+���gQ*%��t_�k�;�Z��\}f﹯�d�����2ɟś�e�����	+��+s�5���	�U�|� �p�ٟ8,YP]��i`sw7���u-��to^.LMI	���l����������P�'|i ��;�?h��o_���㗖��p./o���'̩<�'�6��굍]:.-,!�h}��6g̘���A����ui�Yqb��e1l��;����.�9�������n��?�^�����GW�Ǩ�3�;������R\�L�-�X�.���?��Z�~�#K����
+�w�5A�[���s�b�ѹ������e�TF���Cs�C-��'�F�[E����Ҳ��_}W���ằ:j��*��i�[�Ť�%���|����6=���sd2a�kJ2�u	��(¶rIE)%�=>�;��O��]i���]����׺Ҵs�����m��	O.Υ�z~/Ӡ��SYr�u.�?����9�suN{{UH���G�{y��M�̀3t�^]�/g-�o�9Ñ��h�[�9x�B+�¥>��J[�ku��u����˨q�l�
����oѭ龖$�|���M.NE�)A��\k�՜u]]��R�#��Nt�H���ȸ2?[IW��]3X$||�CD�e��lO��C�y�IE��@{�7a���'t��)�#���*T�#bԟ� 'q_�v
�R���o�p(�#��R"�u?G+��gt��'P�����o�n9��w.�bB��,����?ݵP(n��W����];\E����UOv�=�jL�ŝ5�W�����E�)�M;x/�_���Oy�D�7�W˰f`��y�:\�O:|pw� �s��L~�Z�y�"f$����<~����θ/Oɟ� �{��^wR&��&n�1�g��DQ��?އ8�%�����w��R4����_���0ʄ�N�q��<P?��C7*B�La��]&�7���Z��=��3+ncD�+�2/~��C�����p�7�+�V����}}^Fa�j*t�� ̬����&!�2X�B��G;��q/�U������\ƃ��ˉ�K����ɶ�3�2���a��ʈ��<DU�M��.xn���9I�����i��)
�vگ���k���v�d�{E�%3n��E����%��JJ<>�Z�c��սI8*�s��{� �~Ww2E�B�\^���i'Y�\��L�k��6ٞ�J��g�S�<�۽�z��f �BR�?n=X��dX򈡦%I.��:U=P��@���2д���9�%�C��D�ob$P�$W��q&x���a��rDM���{O��i��y4��r���6���P|s+]l � Ag�ROptvt�z�$w rE��pɥ�ta���%&��bg�?L<ѣ$츢ᕨ���0�R掁������~��ؚ��ռ�o��ٯ�̕���ޒS>�������dB]��h�������t7��Ç7;y��{�i�f+v��w.lxstik����öy����Hx�����Z������Ǐ��1 �y���V�;����8��~!B!��Z�i�X��7,�tO�ۮC������r��Z��2Ȩm?�����r�ps�Lވ�8Y�x{��hG]�D�@����|�'�
���9�955դ9^���c���KRRR3���gb'��[<w�D^_����ZO�o�;n{9I�}0D��D���������M�_lV���u�G�} ;N�&0z���}Λ�+�_hؕ������Epy�F���N��O��8-� I��K�$��ꪫ��w?=��?�����`�pn��kg���ov�k$?�V���?�סП�aE�]�r��ٚ�9-�� �XFg�3Ort��Fdd�l����aFY+��a��JO��{�,�˟<Y
� U��mDք���_��]f�Q;�ɰ�qaO���66(��z��F1G�0#P�Q�9b�79��!$*)+Slm��p�w_��^W�IF��OO��]�|�q_6x�6�L�)잷_�^��U���Pb�|wkZ�O�ٞTztwO#��+���_oy^��L��b��f`]��zo�V
���Fi����d��aP��TjwЉ�2�L�>Q���������C��MV���eB�v%N�"x�槮`�6��Q�51�!��Qg9���m��AQu�y��u�Ľ�ս`��m��P��q��:���0à�'N�˩|k���p�.Nڋ��C��[g��:�mٗ�q*���P�A멮3��F�^km>�2^�6ִ����;�]��bzۉ���wV���o��)V�1�)P|�A:�Yo)/�o�C��U��kP�S��{K�?��~O3gK�pZi[����&ҁֽ��h�%y�޽�������>�|kk��H��?�3�㛶��A�x�{��N�������?��Ν�*]p���:?y��7�:������ֳ�ޗ��?�D��/�[k���w��># ؑehy!�O?�җN1���y[�U��"��2�Y�X��r�|H��{��M�A�|r����d~i�B�]JQ̸�%����b��m��Z���.�X�e,^a^�Ҙy{���O�Y��/Dh��*JN/8=����+�Z�频�9o�����:E� �mF�/=�����~հ�bA�䞧��L����J���]f�q̕�֗�'4�By���n��m�~?�Wj�oM(cE�*����x���A����5��[i�O����1c����ʭ�Q��1�a�v��i��4���p�aS.��÷��ټ B�)��(��ǔ��nJv	ey'�6W�6WT�7{�	�FFLߙ����� ��ļ�:~�k��B������m+3�DOB����e$%�#�%R�w`^��8>/����2?TwWJ+�՟S���SVn.c��0� z6��݌���c� =N&^���Չ�(��!�3/�5�ׁ�>i������O�ś3��6xeԪ����'������ޘ. U����**��0�-y�,ll1^O"L�z����\.��n������ ���1p�̬,���(�?,�t!���\�LiZ�[iA<$ac1U���MS���:NKp}7��re���t᧼��0��ʊKJc�G%��� X�̒��Nk�+��,#�d���l^C7��(M��a"���̐fa��}x���C�1/�wuɕ��@���%�TR&�ccc�r(V)4~I��rs��ByS�24i�bG\r�s�4�9*EW��)�/v&��ǌ6'Դ���3 �H�N�)	28j^Dy��e?V�ɾf���VZ�0ڔ��_Y_h6+j\�pMY1&�	l���aaL���t&�}r���hPRRw���rg"� :� ���m���1#i�7йϕ�J\��K����B9�e蝉}�I!�w��n��r��˗g��4���,����W�ǔfӋ��aU�	^'��$��݄�y���K��%�*��(&�0�����/|��."���̥��7~��zT���V�i��v����L�b�?h&E�Tʏ60i�{�������$�w[KK�9Ȗ|�{�)�����:���x,�-�L�x�:pA}%q������6����1�1񥘖w)����O�u/�!�����"�pUrp�
x�ƨ���?���v[e+'�S�̏���D�c7C�:�?���w+�Z_d�tނ�	���*�}q�һ���>5�ʖWVƆ]K�Z4Iҥ|[t�xK���<�D����
n.镻N�ࣉ�W��i��V)�T	�H�du�aZ�7~Ah�9Xv}}T**�򻁕���d��@��7�4�̔�4W�c��a�׸𡻧'�<�&CMM�>h���BF��K?-]:�w6/BbV� ��qd�����"/$p���	70��:�Y�ٗB�j�:G�;��Q��0���@���7�ď�����vhH�˳�DA��|��i=�,��Y�7e-�$�'���o�^����9��쐀���;t�AN89;��O57�Y�L��x���H:��pY�mF!��ڎqQ�=�5�,�f)T��~����`蹤�1���̀��ŧ�������6�G��:�T�8%)��+���e��,�---UZ�232���f�7 �"m�ي����p.�Crs}�e�BR-5����� `F$dE�ɇ��J��ܠ@+W���J�P� ��h����<a�V��0��S1k��1GH���:� >�)��i6צm(��j���9~$ޤ���!���l���|��_�~���,��b�\l9��~�Gx7ת�N*/�����\J�d$u*��V��W �Z�]���sc-I��C����	�˜�u=(K��:��'�Rܼ�FO�b0��li0.7aR�5�\�T'�a��)�E�4������K�̞��M��l���#dE�,����Oh�DDD�\�	��1�����s�PK�yhJ��&�����ƕ��̦��� Ω������V�$2 N5�J1_��
�"�H	z?�5�zR�f����P��o�v��U.������|��$y*G���k����/]�g�M\����2�l����	G����,vc+�#E��S=��>;����_�����|X����0Na�� ��2��M�k/���_���;U�c�[ǫz���=�Z�P/�܉�ǵj�[����G?��]�����je_-~s�������	HU�L��15@���?�F��O �RȤA��f����K����̂fL�i�G]�@�Jڠ�U�Ӎ[{�@�g�K���qRk}�D���L��TR�~���2�y�??%�_�`k+����g �VC�)�	~�O=�$��L2��g�6�I��t܅��x��F���]ggg���O7�>�p~���+�Ƣ�%rxU�(B^s���8���X�cfgm-�e�ga�����Ds��q�xC,+`��A~^���Ƚ��bi�S���u@�ц�mU�Z�J��jx�ԯ9���
&|̖�0|R��0J� �e�����67i�y�Ns�r�I$�|�TH3�hⴒ����3��B|w%�|-}e,)dDd�C�X
I��v��#��Wi����к��������v{`�Y*84�8�����ec������㮏��8�_7ӹ{7�p}�)++�b҄�r~w�� ���[��R-���P]����r_��u�����j��\	�\	�
w����r����H�c�ۨ��2��JXⲃ|9~۩*����;��1_�Q�0]����pi}I���b�u_	Z�C�pnq�U#�x�C�UR��h*��@��X�&2�����B�y��?b}�6��/���/��v`
nq��>������p�\��3Q���=_�@B������@ ql08�8�i�14tl�1)���s��?��P@ZҪP��ϓԻ2��<��	?�U�$�S��u��KŮ�Q��&ǁ�4�k�ڽ���0 ����V�m��R���W㥰l�i����B8� ���d���9Z�x�m��J�ˇI'�����`���#����m�*
q_!�oe���e����7&��|,9_oN��:n �5�)/D��o6e���Q\�t;(��?�r�{�UZ���۟Q���{��zF��u�#�H��a��ؔSDf i&���$=��UW��L?Ǒ���2����+>xd�B�,PN��_.L,�iP����cR4Ji0&�@��	��/�.�e�1v-�;�V���ճ�j��o��C6כ7���	!0����
�W��#g3��E(m@C�{�������EYdS[��jL�f�D���Q:��
�0O�--m�S�/�c�����]�2�+5R/Q���4yl��J�d�)��bY��l^c3�Q�/�Bʃ ��~���=�z��w�J��N�� �rp����E���\uc�ڋ���y"
_�s��I���&d3hV�B���@_�;�a+++%�o�9�&���9�Z����q��d��ef8�Y��	�I�JW��H�58�se-���}�؝���l�J`�J`�;ɚ�Q��,�b�p ��sQ�y�����.�c-����� 2�g�&%�9/Ĕr:�Nv�a*d7��b*δ[��Vn�W�s1I�-�ׂ�qI������VGb���q��������	`;���%�0N`+�t�N��L�\W�Ҭ;innN�����RNjyX���t��
%�����VR�)? !���-� |�q��Ѻ��M�@�)�"y0)���A�IՓK���C�R�Xm>�'�)o?�����afc��|4�@D�/\���:`Y���Y�ٝV��؍���N��r��Ŕ$@]��+ ��I�_E��py�V�*/�f��s��؝F�y�R�B�ǥ���t.��)l�!@c�����B�/⿘�&�; �&� �cG_��u>3��o������O���Z� ��=�ih(A`�@����:�kU�������J$Ջ�]/�o78`�[4�K�������0)�2j�?}Az��X������3�$��LMO3o���L�]�m�
		ܠ�3����VR]\;�y�����ʀ�{x��%�t��J�2���{�{*�\�ҏ�V��Be����^��5�rv44?�n%˼�*kO*?��8H��j^(p]0-��
��>�u"�E&�Q�s+#.���&���=���i'�9i�@�]\]��@fwtu �b��Z���>�,����]��n�P1t&� �S �=X�\��H��?b�b�G��㳒�g���p�PӉ�)5���I�K�O�Ĥ�on�L3z�����M�~|����Ni��!���nyг.���u4n�߇n1���:��W��7�GHL�G����\v��a��!Prrrj�&�̯d�x�=�<Zש���#���I�D�ۜ�Gq/�j��d& =K��>]��ϒ��J:(-����/;��}�d�*��[�ϐ��l�¦0�䶦�TV�=����n��T��Ӣϟ�n%4 �lliy~�Dj��~3_���e�zX9��ұg�M�V��`�^��� M�h0�����ׯ��M
m-���D "�!
��-�s�J�8]--��6�¿Lo@�|_�z9�h�8���w���o�Mt�9d<�(������F(��	O��E2�6���=d�1L��#Z=��ׯ���	��'m��ǩ�}ț�͑�=��ߟ��'W���*�naD���~�����,ڄ�������ʂ���H:��egg��RHζ�8���)���HT��;m Ē y�/�'��Ԝm�^ȟh�  ���,�ײS����=w��q�x�F+�E�]��l�4��D?���3����@!e�����-���|zzy��'1	Y��P�����;�n��ipVSUN���l��8�>��ͳ���`��y��~�m�53�J6U���-�WŶ�ذ�V�4�� k�,5'H�\u���Fҽ>�� ��W�$���;­U�y�d
�c����p���c���Ebg<�F���v��;��G��P�@�M��P!A�HOu^w!ȿ���5Q��GKA� v�qFw��~�>�va=��4==N�|v�R�4����=��	���%�7�ίF9m�܀����L����6s�s���5Rvhs���0��s*F+FsD�e�.o��,4�����L��L����Wz����ꑑ����Vއ���Ģŏ�dT�e���{��$�Af��JE��$z��^Q�%�auxW����蠤+�;�a�z{�����m�����������ZY[W_%�����x�Z�磸ϐ��ڃ>��s��p'��|�?��߿�@E >^iD�MVN����uq9����/������6(����1�m[k��$!+��W�׋Q��L"N�fq����e��هg� ��r��]��0��]���S/)�a��7��t����h�G��A.1�@���FZZ��$pl���?�2�$�Oog�5���ww2NdT$�х��<�.�������4�i���y��t�
���v�]h�	\�y󏭅H���Y]�A�p%x0$x��#���!��6�.�xIϵ��?Ӝ� i�`
4����s�՘�qO��@�Ij�?���MQ��ޗ5:���K|�d�7�$kYHV�t�q�7 tP
*wz&��J���}]�}�X���M���T�%��ѹ����)�1������I5F�E�3�/c��}�xӦO��|z�ɝ�L�����&ϘƔ�N�0��O�@�1�&Hƭ�T��) �ׅH�1��ԅvʘ@3L@@M{�ݻ§!��ff���lE2�IZ������i��_�ڊ���+�!�t<�;Ԥs%KN8��r�
Z4�n>�*��ֆ,�%����ַ]ls�y@@2jJ�sH-�@Y��E�%�����)�; �s���"7�!�;�!g�����<
�=}"�Z�G�t�Y�y݂GIݟ��o�E0��C��;::� 'cJFϖķ������=��JcO�n� �A�L?�z��n;���}چ;MtqZ� [���[S�3n.�+s���Id�F%1�eђ:����M�d�<a�0��6�	t�4�}�˖}��4�i9����� �&:*���<I��Di$���I�H��Vvtw�ұS=$�T0���u�Jz[@6o�M}ٛzPa=�ĤC�a��=k��H$���d�s��ZyTϘ�Gd�V����r5���+�~ ]�}:�/[���O�l�bY�ģ���G�X�=�e���M��JL���!j�m�����^/A�#��Y�b����A1�w�����6�6��#��q���K�"�- -��3#۲�h�%�vvc��f�9"�ǒ%y�<f�(��@�fg�T�qs�4�lb���g����1㕙�W�ܱ1^ G�����DdT�P��L�&���F��}7��=@J�%�G���4\�96Ɲ�˜y���lk/h��O�ʕ ���o��N�o333?��r(����Jz�g��T����ʣ3ʭ�r������ڊ�٥���J#Cn��y%}"#
DK����Pp�����?I��ʭv	��m��[h�Z��EcC��?5m-�N JI¯�7�ݖ�u!�4,�s�E�xt�0�R
��@�|ݥ+�&:/�� �;�d�ۊ^��%�;�j-����]����Ro��[��T(�}y"�'��t"�}��{*++A��D7��*�����%rmQ�������^k�7C�J���2a�h�H�%*$Yl��:n��M�+ze�9xm2�Ɔ�T���݅������ѥ�����B�����N'㙃���7K�SI�r��c���a_6�M��n��K�>��^]�ƿW���s��xq_q����%q�5 0D��=�?��~�q�j4��m;���(�#;��m�|�.ݽ{Wc�:�o%�?��:"d� ?2os��U�-ζL$^�S�U�
������/�f�x30�K���ޮMj�S���J�"���!�ӊ�@�z1%Cpz��r��?��p�31݄8�@���J�DZ�c�G��Vve���p:<7���[S�cCu����=�ۚA�ȣ���S�&��~V� ����7E��5��O�r񇭕�3R��Kś�������$
;�GL#~+�a"�32;+ |P}WI.ӹ�7��?0����������f8�O����(x��p�m=MTLl��M����3���?k�;We����>�i�&J�^�fT%�^�z�Y��U)I�m�x�Ʃ�ӂJ�wk|��n�3���j�^@�We�yLYn��Pw@�˰bg�ڨ�� ��� ;y��1JѨ�v�[�C��;
�/�`p+E�r
2����Z��/
§��>�#8��d�Y���SCM嘆��?�������/k
��چ�X�u�l&�c�֩e2ET\<hpp0:���<��cAΞ|.j����l����1�ʶ�ķ���ȅ�oS���Lo�x��wB<���[��D>𿆔�g�F]�uw�^�􇎴���Ȱ���8\�Ӊ_�{2��1
�o�� �&�kdD����5�:�蹹�S��9������������6�z����tH����������@n�xeR��kY�M��w�a0�.R�cHy��}��򎀇;Kb����?V�5���=9X<���2����P�:V ��}�m(����w�ɽ�r�&���J�(�du������+���:,(�P@S󘦡>�_�	H�~;�$|��pZ�)$t+ʛȼ��s~�ُ	�:���q�JHC�0�b���� ����F���*ٲ�7��o�6
si����	�|(g � ꡧ�O�g?� )N>�{�)��'<�c# ��e�MI;0�thm!���Bh����X�'�1@��2\8�L�hH���V*�w��..��	>���,�=_��owo΅��{/�}�maA�����n:\�qG&��;[�pLP�e�>���]���o�" ��=�0�J��֪a�P�o�aBQ�i��qa-l`���i|��:7U�r��O��Ĭ��BF��YRO��5�v�
�NH�%M���ځq����v��qߎ��Y�#+6jJ�r���nT��T9�%�����[Ȃ+y(**�S��V���ϟM�m���T����9m`��%Xʅ�`T���� � n���:������3 5*M�g@6C�_
��HE���.wY�<2�=n|ٰfsc�BFh_~���D]��N
LP\½m?*�033�?�8ĥ�b9QJ�+�_R��V4>^j_LK�r"��>5m����2vvv6%��>9��z �Ҵ8��7��c+�v�\�W������I@���]V��)Ny�6s�{�RV?̐���Ve�#�4?��O�٣� >2`�Hl����rϔ�����S��۽�{O�F�Y��m7v��6b�))����XJ���i�����[^/�h㴌���?�M�ފ��r���}�+�l�!D���o�3�(�h��$�|���b�8��"��3�/z���a�P�Cr��I]a��S@��8-�+�A1u/M�V����a�NyHŨ((/ר�
�-�މ	4+(,,��
ݭO��v	XO��2:�J?�~�]��/��^- �vM�n��V���7kz� Sp \�P�#��c^���Vut�����Ɇ���<;�p����˹Y�K{�?�	G_J��m�L�X��j�f����<H����4SG�A'`iS���a��ɊD�X`�Q�ݿ��C�����jc��ذ�|�Ky��9�0�9�Ey ���P�(qPuu@��/ܡ�������n:�N�~�����zi3�g{6nď�Q���D�,�QO�=�	h��V-�1��g���bH|/o�0���QW�\���=��]���JP�і�贊��&�/� $�sr�2�	܇l�i)��`�Y@�	�jD�i3��}&���C�C=���s����)M����W���`�^�E#�P�=�i
�B��r���Hd;[�C 0AƏ�8,�/�h����֣z���h}š+�($s��bl����Dp˜i�=@KK����Sz���6z�3�S�0�Pκ�m�~�[I�]��FŽl��hu~eE�E寒��g�����!��l�ν�H�/�P/�v��[`ER��$*�kF'���W�<��A�u�Ng�&�7uw��Д�E_��i-��8�cRh0Aj���1�8ф[���#�j��N�M.�����Z����sT4�.+H?{u�BlO����U��-N���1=!�������
[ѷL��BGWW�wµ�{B��Y�}ֳ��#��s4 �sG1�� ����7��14��  k�&_d˦N���^jO*�i@����=�:���+ i2O-���By]�MS%�3�+�CC֏q���,�����?M���5��X,�I�{,"��L'�㽗z��aXf$���u@?������ُ=���H��Q�����O^�:������aU�"a���O;�E�d��d�����g�A�@�!`�t�/��>��B+j)C(t&:�u^w��OQ�~'O7�S���̬/�l;�y
�=�8���TH�}b��Rk�?�P{���]E=&eV�{v���N����p�H�\�f|���	��yK�㽋o?'#�ٟ��Vn.#�(D�)"�R>T�h'���Cי=��s_o��
�ޮ�?�S�f��g��yO �lll��F�x�zS���㷇����<�#��������G��Ӥ��V u1q�ۨ� 
'�?��1vр�qp 
C�F-0��*hO����T����u�+�s�S�f3���H���P�u:u���wh�����~M}(�I=&E���V����EYd�o*$_�Ny���j.M��8!ZHdP�(�
n ����[?��u����FS�y��� ��vEP@��MĈ[�_�+?�l�o�ֳG���1�R��Q1o��o�0N�񻴱��2�����=kԏ�ɁJ��m��������!@`��+��v��o�nr���0ۆ:� �|�k���oXh�2�+�a���hG�H�du�EX�Kn�0��e�V�����S�}=_o�w�`�����z^��}��]:<
0k�;]9��s�~���`ȧ�#�����0~L�.uwnɨ��g�a����zT%�3%���G8��r���������?����Y���j�5
�?�����k���r�����;��;{�cd��Տ�[��A��][�z�}5�P�����%j
*�q���_���(�A3r�D���l��p��'t��B���w¼m�\��������ͻ"�h�+p�_��N��o���-�'(dm^d��$q���N��R�a��g�^L��ټ��n�kj���0�F|t��hwK�[�������O�6�m6�m�"D�w���z��u�:�^O�����ީ=;�矟����w���>�+�>�@	��
����B��h'��M�u������M����hgzKQ���ݘ��.h[��HXWs�_�;���(���y�ȩ�c�߹�$���ѧ�W������iJ}y??��5{�f�k��x����5�Nm�Y^l:�6Hz��x��T�c�C���uW�~s����kѺ�u�Lյ�5��0���]㏬�T���X��ŝO�ݝ����W������V��[S˶����1���9�=}O�Rc�x�͍ᚐфg[�˗/��\z_J��y�����~>k�f/��8�a�<?ߛ�^ӷSћ��;p� �9m+5��]��jt'��Y�.������e�m�R��v�֫N#Q��!�����E��nR��f���������@0����C�����=מ�o���8X���૓�5�_��5�_��5�_��o�yʏ�칆����������������x�>�{sH���C[Wk(|ˆ�gj�ѿ���# ���*��g�)4{m�����m�fd%��z9
�T�����ݢ۬�?E{��w3�)4�z?��[����Ƿ�n�y��~��:Ro�QԖ_Vqc��r�"��ջ�}�/X���sU��O�S[�}3H���L�w��uUY�!T�4��������
�O%���2*�7�=�� PK   �sX��G��D [ /   images/6e0c1376-732c-4f61-beca-ab02432631e3.pngD{T���>R+R"H�� R�]"RR�]K�ұ�%�JI��ݹ���� K7�������g�px����;w���;wB?+��>#����+'�Am��)&�,K?�����3
ʇ����Y1�K2i-5{wc'swwwv+;gScsv{'˴rZ�����wo=͌�Xw�٢���!���H�Oo~2����� �� NlE���gp�?}�����1}��o�q���lqwx���Ԭ82�̊!����h��x�e�2���a�Y��HA��I��ۢ/�����cV�폿up�O���o�����a��v��f��J�[A�T:C���c(����N��&�W����
1�2(즔�S�ѱ2����_G���M���C�u�3��v�į����o�-����J��-����%����R�@5�FH�-3��������I(��s^MG�I�w����\|�)�.�'���	'�駾l��Z��tuSr�~�g�7k�Ǟ�������Z�׎�����}�:5�����o,Y�I�PGEEiw��}������ĕ
'�o��������{Q��A�bHa�-��c��z�=���'���t�;�@����d�W�6�S�j3q��@i�.��y�M}���ų������ଋo9�&�	��[��&���p�� %��^}��>;��B<?��ʓƥ���yG-��޼�*D=�T-���ڋ5���މ_D甥+�jgZ�_����nB���&D����T�:���ej��	�Sm��0��tJ�Չ��K��9����~�O?/Z�}�K����z�}=���f�a����A:G������oT�IYdБ�p�&����ؚ^X�˫�������-ر���0L�*)��X�B>Ļ��S�<��?ͼq���e�')rL����a���B����5I�ϻ��&�D��B��N'��[3���uYhde)*+|�{�%�.H�r��d��c��8^[�q���:c���}zY�Vw0�&�X����	U���Z���g*U|
�8�Ӊ��*��i���G�\\p�Nn�v�h9_�δR�6a�5���)v-O��%�w_�`UJ���hnO�g<ē&͆v�7��:I����9�*��\�����c�l@��� 9X
0�Ϻ�clao�Ƒ��-��6�*/��c6}�����(PV<3�@�(��f�v\!u�?+���'Po5I�42����w���#��~ƣޢ��V�h�q�������_g��9���_<�T���+�����V[��]�g٣���W!��ּ�5��9�w�������⸜�Ę��|+���?��o*�Ș׼*e^��6VK����#6N}T�Yu�ƘA�R�Ww]vQ�?���b���.1u>><�y)��Na�qZ<¼&�d�6'��!�]���� :�D?����ҰZ�Nׅ׳��V�� �|=zO�ڂ9�� �2���Z�36S,�c�Ũ�۪̞Ş�������6��Kj
fa�C������)�>�5ep��J��_�ȹHr�Y$�#ȳv�	LڍQZ������RlN�Q�:r?.Wmס��!U�E���Z����V�m t�_�f�M�� *��w�Et������O|����q#}W�}��n��M]�2:8x|d"Z;�y�c��U�|�Ð��v��H�o�K�k��њɷE3�����oOOʩ�d�h�ږW����oϞqPL����$;�W����g��{\g�OV���\��*Z��{t��XFT�y[�fA��n�����-��$ݲ���tg@NgZ�x�������t�x&��"�f�F�l�	0��+���o���D�}އ��p�kR~0B,7�x{�ʤ����S���v_��iLD=�na4�]U�tޜ�Y�:���M3ak����>֠M#����������z�wM<VqY~��+\�P*��pQHxnߓ��-�ɓ2����8�#���F����?h������qت&�}@S� ��(���6��jeq��,����N���S* ��x��k̅�T�zs��SP��w�lt��QO�ѝ�>���� �K�%J������a�n�_gǴ��:b֑O�|N/��Q��W���8[�����5�:�y��u������F`�`��U[�~�&�Yj7�%�o�������(î�}6��P�o�&D�<k)��,⺒J�9�|�e�� d�6��~A�U��H`y�;y�Υ�����oD���r'�g�
���ged�c� ll�=φ�]D��fOϖJ;��m�0�?OW�jf\~m�����w/���X}�7�̧lp�:�_m�j冉����}7צ	��}t�Ù�&cw�r��9�c?9Z�uʯ-� ��ݲ�t������he�-�4D���]��M���m[�ԫܩ���B�]J��o�ס|U3ʒO��u
��y�F��*a�+M�;������"f;ԻU�(�ͽ����R�C������O��^o�u���1�"Op���jD���_	 .�%��"N�Y���`�=�պ���O�ك1��RK�٦�WP�ka,�w[�qZ��/�N]�e1�'FQ���@�pm�.��d���V���?��V��������������?��/��`���fy�܉�����;D+�e��>��2G{��y�K��̋|�����$�a�g�j+ 9�	��)ׅ5{)$iM[�uF��ܣ��!l��	�}�[��X�e�V�'�h������k�y����51A3^*漠�2�,:�#�V��
uQ�k\W}��Zݡ�Ăp��#�x[7Il!�m���e��XE̚�+��Π,l^�^��(���~V!�F�d�K��Dg�+ ��s �T?���m!fZ鍕!^�K�{@��/�v�2�B�:[�Y�\so��^����S�,3~��G0�f�I1���F��s?��Z��TqE�7�&�։��0q�����ցR7r^�U�,+��N�U�f���#B���� � �s9?)]�f��x��]�t�0����գ�rW����}Fxw�&��+I��ϥ%�a�MΣ���_"`���2�C����Kz�����3S��w��[p�Z���Lp�6��Z�e��k��L�ַ���-e,�/�^x��������%�����w��;����;��N	Bf�i�f=H:z4J{����ߐ�A�p1~q9�^���&����8S�-�O���&PC���ED�/l�o��ёІ�TR:��8h�n�{����+@��[�(щ)":e�ȁ�u=W�飡M�S|�Q��0�]W<�����t�a�(Y���=a�X�=}���f�����m�ǐ�Z�g�F̀i�{m�	Ky�*���*zr;��>@o.ő�?��?��o�h9�u^Ills�1�c�6(_�vl
<0�\����2�sE�bF;2 ���z%!>g���Z�]���S����ju|��m�����[Xر�Z@S����u���SW��Z�$�V���u\Z��X���z�\D�$H��壴��c�(�5��_!4�:g���RǬ�Fuկ�C&ii�0|Z$ɽpe��Mm� ��~�z����0�ì*)�\&I�ޯi���q<Gd-��>�c�����p�|�E:gh�g�̗��I�smj	A쀆�8��F��_j#=ӡ�}�J���ޖ�d����������K�[[��M��A�^+=B���n��I���� �읔uځ�;����v��h4��\ �R/�>��]c�(֫�x��E�2�lw�Ū��2
����9��B
�SGqsM�lוq�1��o��6�k5�ʡ��T�3>���E�`m��=��H�]�tF�wvq��ʙ�y#��3���Ƴ����@���AѸH+>���k�Cʙ>���'�A���Шg�h��}y��s}��N�}�袠�;��<�Or�M�병� ��m�PdK��5:�ԡ�=g@RyG���>����{��uQ'(���E�߂���٧�Ş.��	3�>�>���lo`��U�Q�� V���vIC�%���-�оO����]�e�C<�rhdH+��_S�05�CW�X1�����Yo�g���FYo��7>�ôn���z`1-��$M���)��Y����C����wٵ��6MI;�x%�6�\�>DJ�gL�Է�V�D-X�m����K�Ȩ�-XM��P�n�|�\�ˈ�#��"޲oV�q`H��u��#$��v33�<�geE�{m�{�	4���~j��Z-��j���Z���BB�C����4�3+�	B/?!�L2�!�lc�=nw�Ky����` �ϑL�x;�Pmal �Y��Mk��X��*���Fw<��30\e��(|<�>�`��7�`�6t]nV:�+��1����^��
ޚ��U>ho�sm���Mo2D�a��|^egN�Q�f��(&l!��>o{[�;��;� b� h��/ñ�� _����'��43�����gg��ʎ�Qߥ�a!׉[C7$�ɐ��M�P2�5���]{f�Y��O$�a(�nY���V�G�7*�R�$C�w��������-8��d�^�0��>��j�>l���`��'#���wFž�n|T,�"Y�/��\C��]�3���aJ0ɑ�W���m��'�]�|ה�m��́X�B��_K���F���b�����=��u#��`���{�6vhm�|W{�L���듀�����=�<�kX}��������H����Ȫd6�=���b���5eϒ��E�?�Ek�O5��5O|�H�EO�3I��^��!�\1$6·��-[KB;�U���HB,�Iu�t^��1I��Ӑ۽�&��<a�"�/į�1�=U��i�.��¥jZ�F���!Vp�n(��~-b>��P4�/A���iAS[�~o?+y}!�
�O3w~�ڄ�u�Py?|C;|c-�0�[^Q��`?wv60��u�5��=>��&��в�g���r���֡���� ������FK�y}3G���+���G^��,���~���E���͢���������8Ҧ6}T�n��Ș��k�N���l<kZZop�l}zN����`�����|�ӯn�I�u��g��}� �٬^-���c���`v��R�'g\+RB�J~���nm�����;��d�`|3��7�R5�x*���� ])�5��w�_�����/;�k9�Lb��Jv	�(�7q�cgڶ�D�4��#��Ge�޳S��d5����#���_.9�HW�$��(|z�\K6_�7�_���J�|3�<��k��iZ�x�9��/��Ѹ\㎺���MK1�
n�����~{,C����'�	iN��rg��X���6�}z��z#2hO֌QЉ�>�<��0xkԘV�ЧX�,ߗ-/�F=u��9�'���`�X˩�ұS�v�G�i���V����Pd>p	�Mn2!��Юlfl*f���X�U�p��9�\��j{�lFf�~�&�C�#��;*��Hj�F���>��6�&�1~�.{*�_��RmE�]O�rqYI��c[e��ϣ�H�^��5���I���;��T��{B@_o�w1s)��{���}7h&v܊�>Z�́���n��ɲ����O����{��QluO�)0�D�:��J���1�յ��QZQޠ�?fN���#���lA5?̜�&8#���-"�����,b�K����>����I�"�Ӝ��l3�fQf��������7���u����R��J�.����5�60(���>�$B}bR�A�7�<9!��x#R�5&~{#�n$L�aq	��"�(���t��R=L�K�_>�p�����V�q���C�pPӶsr������&��'B8��#���l�Uf^ݽV��C�eC?��(%�t�(�g�v�Z4��U�@2��o��I;s�;;����������#�-���{p�� ΪVsV�RvA��T���W��|�H9M�S�*��H�#�yU���p���8�(i�Ju9�OE[_�\�
�ů��0��Zr*�]�/ �.��h����^��&Ź��;�f���b.�V�E]�U�up�r{g�d��|�7�������ʾwO�j��L�^��f�K�5v�����U�<W�����q����B��1�����R�������[�%d��R��_�TS��)�:�]-���gzV;9m����iL�"3������\\�+[����Ѩ\	�4�-�/5u��Z���-�=�V#%J�$��l��_g��C��b�����pǔ�8�����x�&��P�gc2���A����~�%�ٚ&����\+|,��S��Ohf�=�d@�����0Qvt�	,Ȟ������OG��R�:\O��~����ҋi�Vg=`�����X�����՞Կ`c�5J�����w�����w����Ov���R9����Ǒ����͘�L!U�����m���w6tHХQ��8M1��d��̻�'��k0�<5bfyaE�b���煶;�&��� y��W����+�1Q�GWGW�]bKk=�u�>�9M���UlBM!���#@��]�<��W�G&9(>��٤������:��%�&}�f�^�����������΍]�u��Z��D���?����wG<C]�ѵ�_{J��V8U7�çR5�ơ��L� �0�G��`����
׍F!���o�g��r��_�=��3�؍J�d����m��VW嵪 e�x����/��C�I%P��!6��H2�&jr�ܾT�?��u�~�i�NOX�>)����4�	�6�ݯ��AlmWZ�y�p|��xT��Cf=����w˛
���^� o�R̓Nݨ5σ��N����=�JL~f�m�MY����ӓk�y9�V�."�W'�g�5ro&I�GMa�T)�{���D{�k�p���P������F�w��,�[�{��#"����8��;$����8�y��L|��%�`��C��Wױ,uYň��g�6�O[ ���AƑ��͌G�峺�������c&s���[�ri 	ˤ��D�K������3��`��_��T^`�q���:�s+�G�"ڿr>�SGv8�F~uz#A#w�UTw��|;߸���d��K(��q���(�k���t}�k�������)��Q|��.�� ��ƤN�C�x~����Inyc����5�1l��B�C�D���.蚶��~r-���}���ƊL3#0H��Dob�a��t_	r�)�4��n������x����Y���X�q��_���H#g"�^��S{	Z���D��]7�fd8,����R��!%&�zS��zڰ���^������+�i���q~�	$�'��+�����L�JQ��/��ylu,��X��Y�3�'�_��q_6��\[�գ��zdԧ��7gR��T��5
�T5vLѠJ��C{��b�i���&1�+���ى=�ϻg���Z�Y��ޟ��G�9�]���1�|="�!�0y�,@�h6�"b��!Y��7ހ�ܻ��ė�(W��~wZ�FW�ƃ
��'�ML�!_���n.��h=��o�ܑ����!�����-�RQO?��1�D��3�ch�;\��YNb��vt�r.�@(*��^}�p��_z^#Qa(��j��a���+2$��3ө�ّR&�Y,@:�q�Ӂ⶗oԙ�i�-�K���?uQ�������M�i��|Q;��M�ɉE{�Z��k/��'�O�	x��(>E�w�D�!k�4��y(.��ޛ���.&���=3�7[՚k,ijqq���$��i��*0�^f�Zw�vDG ��~_�r$���2�p�E�N�����*���h ��,�����msk�_;,l7�l���^�[�G��=懳2B���w~F�T�n�E܀Y�c��RF ���Ǎ<S$��!r��Z	S�>�o�4該�o.M� �z��j�j�Dtq?8��aѵ�3�S?�]�Dc+Iw���erw�{<{Fw�v��޷�G"���o%Ee�4����޶�����.i�/Cé������U�f�QT�����q����`��P�D?�{��hݲIQ2&�cD)�=ѱ����� i8mA$޴�s��{t��v-�C5�F�8q�6l�����9/�뗶�b��YP���l4��,��u�Q��J�Zq�?�%��]_�i�~�F��Uip���7BϷr:9ӕU��4��x�mVF:�"ሥ `wk�u�����E��Gñg�����6^�x*�u��EY���j��8�(� �X�𒌅st�+�~�e����:V�6���I�_=�e�X�R\�(Ӑ�
 *XË�0�|6s���'!R����{7T�8E���a�!��l~����9�����6���F�ve�^��9�]�i}�����S�����˦�J�%�/ɩ2�ow~�Wo�ѿʺ�[���)��NI�*�4��:Xa��P���7���Z�����*���h��,���� ׹������_���bL*�'5m�x����<��A��� �M�4�'X�����4[�|$�0����do�j��� ʖ�y�Wrk��X��0�}�v��p�&�}�F����bU�ɞz��]��>���?���� 5��6#+Z��Q#�_�Nj�p�!�%}�= �l>~K��S*��_����鵸����w3�Ɋ��:�^�*sf?3�`ɍ��5ü�6���rK���h��-;	�|�4��>&�hdW�9��UX>����k�L����l�$�Pe*g�mf�kk�(��Ƒ��EP�,�+�VWW?�<�C���7�z:�+92��,�RD���ȹ���\� �cSܛ_���kY�Ok�!�e��'a(_��rrK��R�+��%�v9R�K�_�����bf�7�!�:���D��qM�1�7�c�D�>�)�ks��?���'��C��3���ZR^'���ܕ�P�j]�a�!��T��E$�Oh�"�;`��j��;�w�~����ð-�m�p�4��I(w�r��z�������+��Ƴ}���x����%Z��f)?!����p��i��
����T�_,8};_qk�:��z�T�5l����s�����P�7��ޫ�;���8Sx��;�`M���մ��M�/z�k��):Z�~�Q��̜�W�;�#my��z���&=AYҎ8�xlzq ^�p������Ç�ى~��I�3� ����܂<���w+>�hC�P�IJ���Lz �Q!�
��1�m�rk��k���.g�ৈ�S45���\"qW�S%n.7NÅ�_om.x=t�O�9��B>�$����Yln��l�zK}w�t���S&�Wqí���8�Ԕӊ��I
;j��Oh6�n�����NQff\���������^+���4}���Da��|�ƀC�\VC�h$�L�Ň��]{��@>���u�3]�B&��|�ٟ�I��B/�r�s��Ϭ���dw�.p�~��:Br�T���_���L�Y,��0�	mKm������ipG-r8����'�]ϕ��t� m 'mE���
+2���S�dW6��(%�X9���Gr8}�f-@�\�k�
ZN/��H�6&�͙Ӝ��)^��xL:+ J�஑e����Ǌ/8_��,4�G���;��ۓ��Zů4�q�{�8�3���8^'�ոK_�x�~�]<�g�Q?ղ��3�dX7��'���7%Oq�~�ip�X��7Kh)�:�<�e�l̼W.4���0)�+��!�t[?�p�	��}��R�	���3JhF��a��D�_�j�܆�;�W��$�땿��6Җ�F��P�9�1i�A���YJ4(�&ۣ�4���xHrü�po��,���\T^�P?����>�m��cs�.��e��E�4��==Y�&�I����[73_>����ax��+د����ގ�ٝ��ҍ��{�z�6���)"��2��;$Kd�U�ig�Gx�η_4��lGq�}|�\.W�A�ѩ9��[�j�|u/��^TXu�M/,�L�!G�4��;���kU^��5�6t�5�X�b�l�Ǯ��&�#tW���_(bBC�FR�n�I���z�G��r��������R�kC�.�d�͏���C}�ԆY�{:�@��^x����}�4��(�-�h�'����t�<�����.���)�t<K�c���q��qRM�I:֊��NꞠv\��!��PM��|���^?�5�̗{������k�`��.1�������d�N��y������#[��A&+�X�ێ%z1�_�Y��j�t���YLo�[�<Y=Mz</[�lf��j�q���������j�~�ۭ�w�`��i�[�C<�r�DL�Ӛ�}��_�~k��$�j����Cؾ�ǀ�c���vu��������v��{�%ț�����0[��t��0���~�O�b�HL4΢�nض>�ę�yE����m�(�����$�,��a���˨2�;����W��C^K���	��48�P��ZT䯳ߛ]�����<�^�>v��XV�c���b��.��:��;��l�)���К����Th�9ϣZ0|��8�,�WF3bN�N���]�{�8W��|�`A� (�S��M��m��"�l2� X��nygz�v�`&7����j2��[?)��0���HZ�,�k�Un��q�y��ʶ����aڛ�h���Y����BSJ�tBY�������g�ܳ���*�d�aR�����ܠ\�1�4n��,e�Yoͩ`ӊ���K5m��!�{��N>	�����^�'q�]7����2ֿ�?2�~���=x��
=hp��� �Ύ�/R�S��6�}eܲ_~ʽ%w�����3]��ڡ̘��5n[�%�D��a&�Z���pd��~�a��`�b�U�E���8+X��ݒ�$��>ئ���X6��9�˙�_	��I���O|E��F��r?sO����Ir|�t�T2;׭�4كD�S>��'�����O� �,�!Cv��%�J�h�X>�5D�Y��	����Z�W��m��1���8�������R�������b�u���kj��*X�!���[#��A�V�����(�|o���O�~NN���*�β��o��Q��FK�븎۩�.r�S���P��^�59��SR��}���%��{��Q�6�ש�Ȏ����2e�'�8C\�({���z �vp�Up��Iݲj��UF����絷�J��_I`��e���]u����H��б�.��Ę8�c[c<V���Υ;_q��3�ER��l�*�j�BjV&Ѩ�o���_~� Y�0a	S=b(�@o1����
�l�q�;F"�~M��PMfʂޯ--x��<Vh�2>��kL���B�U������{Ҩ ��:���"��I���R`L�v-쇒��/(�`���C�E��F_MT�n6��b���Z��w��;�0��[�RFw�~�����h�vu���9 ���ch#�O��Ԟi���N���Y]�@��S7��>��gY��l�']���ٸ���[�����bS�OJ�X������EMqi7!M�֨�a�G���x�^Q��T�¯�9�7>
�����U��p=k/E�7��?�d�U�=�Ʀ��"p΍�Q����N/�8�/d���ҊTҹ���H�e��|엾�	l v^����"B� $i ����8+�MJ�	 ��/Xj$����6�9ˀ̧��T��\�2�ػ�w����D�Ч21ٴ����ȉ����0h��l:65��e��{�
��z �d�O�X��*W���D�.��d�[�ʕ6P�ų�]�jkf;�%���㷙~G���n��ͯ`	�`\�O[�inן���^�'e��>�n��>�#dMAne��<�Zv�UR��MH/����P��6�]j����1�=y4��r��� <J{\[�/4f��&���n�;ߡ�.f�i��i��x���q��}��]�pI��?:�Ӭp����q�m+5���p/�x��R��0	��m�F�.�Q�p7��%���L��� 	�t&o���R�LF:��C�!pR�4J�<Q`���,��hW��E��-��+��6jp���>!M�r}7�焄C%�A�o}}�׎2ɪtbx�^iVށ�7l�����.B�ò]�Q?++���8]�~�'�|��/���x���ؙB����b��/��-�GZڼ���F%�[�^>nyhu���}l>:*.�ƽm��^����;�7cqK'n�\L����y�*"ޱQ�h0a�����I
�iY��Y���F�8.��م�ÁKM�}A�|��x 4�ȝ�[�H�qDf�Z;���9��>����|%�
Q���O}��?�0XQ����A����R�x�1?V������þ�ߠ�y�{o��I��]�x.¬ª�oH��s+5'���������B��c|���6�>b�	��g�s����73���dŤ��
�7���rM����;6��u��dd����QU�2`����%%E??��쉻}h��>E��o�t��큨�����~?=&��do��Y$1��"�jHg�_���||����ځ!M/���� �VW�e��4g�֚
�zӤx�!��O}ϲf����;��;����Q��5؞��1�]eK��4 {�jnȋ��/'ؕk_q011Jf66If����/L�	fGR���y��q�LP�qe.�D�
����$wm�Rj�_�����0D����7A#Z׻��V
�ZW�۽  �C�ZT�2P�����_�l����&r[i�M����q��Ez�f�
��j���n��S]�d�}WFSZ�ɉR��=.�x[w_���
V��^����wԫ�+1�V_3��������m����ӈƨ�[����$ ���Z~\�E�O�C�C+T0�숑qz�7o�Gv������o�B�wR�hJ0�%C�ж�N?[n��xU��/�|�3���;��L��M_mI���u˥�0��ؼAK�g��G�O���iD������ӎ	����=��Id랶��6G!U��<�a�K�������0�7�-��xD�ߘ��/����y_!��. Cr#2�ɵ3�2.�IS�p���@�7��0�����d��`yx�2�A*� 6^���j]��b��f(g���%e���)�t�K7��<�K���CO�^�1�#�,�~#�١m�T�1��N}�$U+���YHf��ѧ�il�H��$ԉ��}ڌ%�"��_�b��I�A��C�����no�z�.�%���3AdD��CoqYax�5����{���ُ��))xT�;;��lr;�}�k(\`��p��̋���%�p�3%y��=��etL�������B�M#��c�HdK��H*�i�
^�z9��˄�+��`l�8�Z�`F�UO�/���R���T�r�7��MFr������hǚy�k%��W&��V
:w6>�)R1��i*ˤ���X;��)|��PWė��ޥ�Z�o.�	�H�hWM�J;1
v��,<5�0�YT�T��^o=�A������D<������܈T��~�b0�BXp�$�@�=����yy�����G�o2� Ã�2D�:�&�,����[oO�/m�mRZ��_��4R�u�����#��\<�(�&g:F��l�����'{\���P��5���̓�ٰ���C��0/-xIP�*���#�W����!���I3�|��HV}�h�Y��i	�v_0wa�kT����P��I����
�����/�6��F�D�����OU��X�����G�����K��M�S�	o�7��#Yl����>�1��5O�h�1�l�d�@D��j���j3�4!��s|��7�0E��_��S������ �.lg���f������Y�m��R���[�c�j��NC�Ϸ6;o��׃4/;0z��#Uv�r���K��>��V��o��w�)�K����w�GW|���z���Zn��t�� ������;A)��݄k\�{玐_	hL�VV�);�>}w�,a�Nr>ŷ (MO�q��k�5*�NQ��Wm�/�O*&��{;)$n�al�w8�����3��Q�/|�V��j����<�OeݴG����n�����\/O��-�.)Lx�˷�sħ[�4�S\V�d�0O{�N���P��n�*��ݺ���隧��Ւ��.5�
�����)���j��h*�����a�Y�K�K�
�&��>�=R�0؊�~�����-]��;
�I|±%�{77��?>J⍭ф��	U��M���:����y�M�+���
B�H�s���~�-�\	���=�5��PD�Yu��k�m�iw�5W(�q�� )�D��t���	d��q��؛����D����?r[��}�~U%�U@BS�7�TI��I�Tɲ��!j�����8��	UNA�E]� -�ƎBZA�G��v/w�%����C�j����k�cZ�/��)�#lQ]�Mm0�&�D�6��L��Ը�������b� ��!�x3@�g�ו�Tb�f��!�R����UH��wIYޯ��$8T^�b�Dڨ��VD�ٟg�\v���X�k�!����'��O���k5 ��"�Ъ��.�<�b�l��)����F�ܓv�Z�e=�PYVnÍ����ˁQ�)aģ�.�u�z!R�@xvH=�O:�6��ϕP"{��J�H�$�f��<�����4:i�u�P��羾�Qux���]��W�/� ��ikp�1D/����4��� Mm":!���X"�����ꚠ/ƙ��(�f�߲HQ���v�q׃'V=m�81)���zm$�1��wg<��_�^>�h��N�b~�X��4�7��OG����T^�6O2M[=)cIv�Y�nC�bk����旞ݐ�S��	!��M��P$E
~Ч�1�+�]i�����c�F �$�ծ����ǟ��8Z���C.��h�ط�;u}yRx�n����+!"��1E�/�Z��xS��|/o;~>���tF�j?FW��{�o����v�G���39�,�)��	hS_�ϵ�V)Bދi�w�2�D�IV���������k��@V^���e��2��(I�§���R *~wy���C�X��j[�۷S��~�1÷��%r��lt2O��C�ɤ��J�7��{Kќx{�X�J�흙e�~r�|�v�G^OU�j�nK�x�>0>�Ӟ�TgQBJbn7"��!8i�P4B�aUM7�Z��ee���'��
W�~��=���3����>踖4���A���c!2C�pSu�4Uz���n�f�tuNgZ��}����#_ ��\E@�{G��I܇��;M+Kx����i�@�֖N��3�gk��֮}��(�׾������5��#���;L0SgS�%��O�ʞT����8��Fzܿ\zX��̃��|�{6<�s �zt���
~RW�v@�al���T/ba9ЁP������ʱg���Jb���+�B���o�^�/~0UH��&xa��J&?9
7�w$ב/c(Ѳğ�I�6�u,x�{_��3��1�y�4>��j�K�4��u^��\�k^ʺ`BT(�%B��4��yu���5�+��;f��Q���/�{�K����A�)���_N���0�~�}pt�]�$�7T�?2�]�Ⱦ����fP���4�>�z�(����~��{�4�!X�n�3�F����g�W#�4��}��cD��F���>r�2�Oo�>O��Z��n�W�@Vl�����~3H^H��K�_�HA�jt�|�l_*�����T���OJ���fX�·;% 񌬋iP�\U�q�2t�����KM�W����)/��g�Ƽ�-�<�ix��B���Dp���r%� ԭ8bZOATx�2�Pej�cu���`���̺��Bڒ>.��5���7ȝ����.��N\ȟnR�DE5`�b!u\x�*.�\>.�[=��w�Ɍ>��6�&`O1��IZ}�Q���� ��؅�@:`I]���I��������W3�3<q�nB�z>��*J�ٹ��Z�,�EV���c\`I�@�V
Qw���j������A�� w��) ��V^��)NUW�qW�3�׺�K)6)������W2i�0��841U3� CI����1�b�F ފ�g�o�NP�z0�0\t�D������l�-����[	(@���ZwG�r����|���y�����F10�ɑlo�o�x������{�����ix���T�g��M HB�EH'
WZ�k�I���A4��P����+U�+�+D�K��U��5�sY���3U2n�B�]�+�Enl�a�=��%C��!�����$�!H�}��@F�u�i�i]Y�^����X�>y����}}�f^��01B�f`�����L�h�dko/���-�m6?եa�6�2�>z�Cͻ�8H����n�x������΋�z)��;�̪���l X^�����
��R\�I9�4䱈
+Ҋ\��Ͼ{��>��o���6C�B���$�3v���s-A�ꗥ�S2~b,����t�ƶ|��[J���?����X�#k~0���۹�d�/����-�(��Bۚ�������0��T�
ޢ��X�s^�V��q5����R��9�Q)�`���H���H��׀��e�W���Q�b{�e�à|
'S46�����G�[F�.]��� �Bp.��	N�����=@pwww����� �;\r�y�����ӵ�l�~���Ϧv~�|�� ��[�_R/&|��������w^ˊ���A���(�4ܧʈ�F7exg�\�"W�ށ�)OI��T��{�6H^��띛�A�vi�U�*���d�����'P6o���A���EU�C���f�7��x ��Ԭ�~��	+�fvP�۰K{~h�}����"Sy��ߺ����?e�0��"��ՑK�	1�~0clF�I�XJ��%����?,by������h�f߭��=��DHYt��c(�(/l�Ξ��C��qKJ̒Q4�{�ﾊ�/�z��l��"�=�FL��)��Dn#��8T�	R�KeU��)d%�(��J�����r�ݦ��y���$���,��%9pQ�݃0='CB��0���y�%���x���D�-W?��C�=�$n�'{����e7!��bS>�� �������(~��+��PD}�*�H,B���kS�~a�����Rx7p�P��'Q.��5eJ�E8/�ٍ�]PQ��r�~WWX�1ijiY2?�.���86�-l �k�ƕ���q�����W����j�s8YЌE:�;?�<���sE���\���`TT�+7��c7֯X���ɤA��ա�1�+�{7�Y����)|c-
��;�aM������B�~q!��/���HfH����*:�9�ai�����F�������qJb�j�Bl���b~�Lܺ93[X~-[[��U�Wl_�G"��M�H�,�c�-�Ĥ��;����L��W�yn���C�'�_O�9��QH��[HwB�_4*R�~8O*]�	��ύ�+�-�#W=Yv�\ܲ~�sG�����Λ�\C���<�7zCNY���<I��7.d׿-��cG����c<��-�ACE�+z�pȮդq�n���|f�,j�!t��.>Yo�� ��
�Gt�(pFf�r21����l����K8�~�at\u�]�[�Lplڿ��Ǜrf.�����T��v�8�խ7}5aM�W[�����ROim���Cz�����m��+YږQ$�q;3�lK�����9�
(��q�M �����#|�X��VY%�µ����S�4��L��T�_���\�>)*��	��J��2bS�3��m^J1i�ubYJ��46�y�}�̃���f���uK�*a]�m�����	�ױ1��h�q�o����<u�O��[	�ϵZKzC�FG�Nվ�*����� ׼�RWKHI�ѵiZ���G=��_��z%��y����쐦+ ��G/˄P��(�m��J�:���3��2+o����v�.��e�O�IP�Z"����������5Q��H��D��~~��U �PQ&��*F
��/Mzܮ	X�`PH���������@�p�b�,~$c�i��&�Y�LXRĭ�T�2�z<�֙��U_E-��3R�ח_���׍p��!D�W�Ό�{�<�^>��D�s�*5^G>��d�b�O�e/�p�Z�V6�y0X�jx�}#G�������vSɔ�<w3�6�65�`l=>�kd:�[g����ԭ��vϨ���֯�o��*æ�֛ܩ��ܘ��$�&?@����II=��\F��q3s�m�y��l�z\�X`������1&�讜%�h�}錝��u��'%�؈��ή��&XK+��^ef�����q������b��f���N��"��cJ�dFi����L�
��)����>ۥ4�Ԃ�Ӄ��v�w��͞v�,��R���|��磯ϊyO���E��aO��N��d���U�5|��:�t��L����
7��;�����g���w����ĺ5	�!�y�GT�]���䓓�3��!t����������u:Al��h����c�C�_���ĜL�����K�1t1�RφS�\?5taQױ��,*5�Ë�������0|�sD#M�)�8�t �����_�ԧ�2:j�t����ɼ���Χ8��/��B��,�y�CV�p�U@C-��ն�U�o[��?@<�M�D�����$�:�ߓk�'�?�M�Фp���fB��ڇG�'���Ҿ��$nc��W��I�:��'$i�*�d��$p�X��0�>H�%!�X,�wS�d�b�h�.^WS��E�M��Dui\��^�3p�"�o�������Xb��8c��p1��x���dkk���I���
��ޣ�u��\� Q�p��=k�A\�����©��V�F�j}����l]q�/ީ�ʭm��
��W��F�����_	���-�n~�3)`�V^~�3�sO���49M�4}��z҈䍝��.�frޡl���L�7����?5� �[ ��������['�8Z<�\����VV��ۍ�N3b�{�8��҇�E-�_�U�K��-Y�w�`n�Ҧ˃�q�����]�[���o����T��V�������\B���J*�j&�����V�^~QC�l��v�u���P�y������_�	m[Z6R�R�w9�Q�w����`�c���5�^�)�=EB�#,n��;�
r���ۗ�Sp�w�§[��nʪ(TãN{�d֤�\X����L���*R�`�nC��̑؜�`QFZ���9�]L�k��{��ʅ�<�x�]'r�]��>M���ڬ��R^�:�<���93>�,�'D3?�܆��^���PT����)xL�\�n?����~��>���%5���C�dz�ʏ�'t��anK;<������^��&7g����-|�[�y�W�͚����&���ҍ��ե%� ���=�k2�t�=����>�d�g����C��}��Ly:B�����l''Q�c�f���kQ�����d��&�z3S7kE����]�u��y��B��?�V���|Gny���g�<%Ba���jK|x�(�����!��z�ԨX\P��5��՝i��,���] &A������pJm�b��.�*��|��c����8!�炈1Pj2�#���
l�Gq��cG�ð�r&�!����**sC�DN��^EW�
Zҧ����ُ�R��i��B���Z�뵬���+�L�e s#t�b���0z�B����[JT�n:=�{-m�?�i(�h��-�D<L�9�]o�sAE[� ����|ʧ�M�4�$���ׁ'$ξ�d���>=�<�B��&�M_>�܃z�]K���� �=ϝ��l����j�OhC1oB� uz�,�{�eN�ש�_�j��*���%�mʹ[�d�x�P,ah���T�qk��`��Tݣ٘r��ފ9u.�T��Bx
pU�k��������Z�����������F��ݒ���/ps���0���ȭ���sp�97֏���é��Z>أ��$b���J����Gr���D���T�'�U����y�NG�h{AO��43 &�C$1ㆵ�QD�]Fa�tX�Iia;� YNgoAh\y@Cpr�i���-��P���A�kǧ�ω��6hs��&}�*i������)�9(��~��p`)3�����KĻ�xīZL�X���2���S��hC3o\Ғ�F�Tݫ��È]�����s��u$�pr���W��el��w�~����/qcbW6ޤ熴���b��Y9�P��A�;�]ܻ� &�g<Һ�x�+������q~�ϧC*XB5p������}�aa��	���za��K=��Q���M/�S����A7Dܗ��ρ&�9%�R�ɯ��o#v��KӲz�_��7�{Z�����򻝚�ּص��go�i)�y}}������$$�2�a�#�0FR��:����Kkk{�e]��k��E�!��'�lC��l�F:�f-�q>���.�B.3�8�0,�!���lC�X�jkj���-�E��8Ju��]$��b��<�,ư��~8rF)]�GuZ���,��mF�����kS�q �c!l�2�FC��ng�˔k������p[��ũ�95=������S��O�"��M�t�w����[E?D۱�HE�
Eaظ�
���Y�}�>�R4mX8����a�����_6�L�/c83=��.H3I<4:|^�?��}2ՆB��JU�{�l;���B>��:1�J�0�����g�c��>_�ް��c�~9s��$�c�4�����poI���/���&2I����k �C������?A/�*g��H��F�uZ󕭬��?H�W�R��=��B�?A����D�_r�n�qwX��n ��؆�ks�㻉~�1�Y���
��|�V��*�Z�[�����^A����X���W/�N�~k5/]���x����+��f�������aظ�􏾽FDͮBM7t�[���QP���-�+#�������5��$D�g����w�"�A�OJYFF����{ޒ�#�`����_�7��9Z0�����,�h��vA�Ps�����%�y~��=�}����*�FU:�������7�' �fA� j��~ӄ��x���w���q���gB�o�sR����[���V�MiA÷(�Ȣ��D�M�a�T۳� ����lVE�֠Y��ї�O(�x��7�����/�`���1���>�ux��\d��W�N��G�l��2�O��ߘJ��.�i%o�%���wކ�,�u[�ƖQ�,Wx�AC[23D��� ���e����pkڟ��eм=||���(F�Ӄ؈^9c:������T]��<���� ���m>�
=���[�A��'+��I�7~>�_�by��K�OL��Sf��	m�ES63[@����߁��*/bD9�Õ-%� RFh��߆��!���5ĲR�F����=��3� AH���E�h¿������$�b�{��ɠ��6�9fQ��h#�@	��*�Cx�������<.��=i�^
4��05��:���<QJ'P�3����Uk.#���6k��������z��,��̿|�����>�f�a=�_��U�0�$�r7-�{*Op���[���v!홸zD��z;�Bv�w���ہ�w͢�AJC��-g�2<���R�XR<��#l|��ѓ�@�pq/�	��:q`�B�\y��?�2�uO�᳓'��PaQ:	V�|�d!<#����_�6�����{{��s�9@h~��^���T��7�hQ7����;0fV�������q�F4�~b�N�B��Z��v_��;���&>�J�ۤ0q+��nt�d���$�U�o�q���mb,|z�6M�	��^#�o ra���9�k��%�U�v�Z�px\2��w����aN�,��[���)ė�v*���!��t��a�u2�~���nn�6���������A�܁��a݊X%:�>�k: ܚ}ؕ�|��׬U��:D������+�m�瞂����2E���Lkukqqh��O�����Ę��xP3�+�o��f8��ـ����;]�����,+������2���\��d"��h��ĩ�Q~~�=�㐑�<(NWEN7�TJRj+]���c����'����4�]�>�����g�;1���Ӆٍ_j�x|�{����?+��w�X/
���FX��+擕@�_��Q��oq���W�����z�aѓ�G�%ģLz�f��ãb��x�̍����ٖ-��e��My��5D�@�-.D-�F������
�UQ]<�=����Y|VH"��,�:��:�<݌ �#6�z�Ȥ֌���gn�Z�3*�o���M[�]G=I��	�}# ��v:�4��aUA�0܇�扴Ί�j�j��5�i�!N(���6��$7���l�����n({
�c.�_��{N&cL�&61��Gژl�Qġfr�3h����{���Uϗr~�X ���Ա6+Y���)����'<��/����	�}�%����!:�9�����,]�+>�l�ܫ��qM�=��V�Td��
�Vf_�},����w��WNɒ�w橀΍�Cr��kF09����+��yXD� y�Y���zC��*H%��"�?�	rRۍ��j�5̋4sYɤwE�J�e6����Dr��
��'���w�w����q������8��58p���t("���Gah]�����SK��^�aԖQ<@}d���<01�T��e�������B�M�b����z#k��Dh��q����{-'8
T}���û�Ip�b	mS�F�Q����U>���;���2*�nED��I.:��a��=�ue�o���
��ѷ'^��x����N�3Ji�C9_��<�-g�WسV�܆��~�;0� �&���M#�R I`����bp�9����7��=�#^++����S��;���Ov�%BzF{OO(�}�7�ܪ�I���R�otM��fh*� ��_�U	�����2cN�0k�d�b�)}��Ym5��qh�WϏ��a9���<
޾L����B�GQ/5c�j��&���?-� ޽���^*�1�f�g�����_s�lBR���������;yr������u!(SWޘO8��י�nb�K���q���]_^X�Dh��J
o�8d��g�^��=톙�%�ʢ0z�ۍu�_ҧ��K�u��h0��u_Uwa ���˴bH挶6Se�J=Y�#F)m�V��u�U� ;�7ӠS���{�P��{{�B,��1����:��2Y�m*fi�w��K7��'�qRu�3�o1Q�s��(g�0�߄v7e&2y!�<�$�Qa	X�b'Č��˝�Fᙿ�8�2����E^��U!/G�t�ߗƿC����/�cQbq�~�u��#�జ��Sߏ�qz�x�;K0�[#,4ܽ����f#��}��	��}�Ƨv7�������f�/E��Ɋ���r�#�ߞv�;���o%Mq��WbZ�4pa|,w�,NY��{�Fxo����!�o68UY%���!��ϗ��� H
�]�G���á������l�e�j�>'�v�NX�x� >u�^Z-ɧ� �q7�����Yf�3�ީ��O��\db��!�F��U��v�u��:V�.��=\�0�h���@c�C�e�\��m��r|�+�������ٛ�"�W�~�@;6�����V�hg̃'N��R���1�mY�f9��:%�I$V;&�������.�{��w^ȱط4\s���\ZFl�Z��e��\V:���E��u���:�N
�1�������)��le��:H���"B����{JAe�3=���g�0���"p�!s?�컖���۾���
����	iCJH��������bt�����Q�o��־A�Q����YyϺ���u�<��Rˮ�� B��5[o�6����<Y�/؅���CRO5i-��e#�S6'�]�`��q�����U���}���w�w�]G��?{�)EAՄ�T��TA�r��U�5�����G"�g��vɼ�Ȱ
�� �k7]�s,b	�{��lt �؇�X�^�-)�����B$�E]�XSw6*N��~�0��]F�ý�0��E���D��"ԕ&*eH�|S���8a�,�S=���R4B�����6_��@;�>��Ѳ	�$ؿ�a�GwW��ވ��n������\U� a�1P���@����F�Ԟ���A		d$��ʂ�-CO�M�@���b鼩h�r:���
`ي�]0���N�5T?j?^�!u�XcƑRB\b�)��/X�u��u?L
Y�j8^�#����1	���\�*{�MK�	��M�����=���[�L㉇�B��#��ҫL&��[6�n�柂�lc>m{W��9ָ%�2b�ľ��U�*�7Û:;'����tm+~��� -��]^�P��������/��Y���H�ͻ�;��l��94��'�Xld+��,���C�g���n���rH`q�d�"�sQ�LOt��is�|�&7���v����A�y��J����f��������>觴�_#ܠo�rR��PW+da�����y����i�\0.dh�����4���9��{/�ܽ�f�!�&��zxl��b҇q�0�y~݌��)��T��h�v�iњe'Ś��Kʠ>�] ���Q�{������H�%��EO�lۏ�����0�&p��G��aLȥs��"/O��|@EA���s�����L��T�N� '�EOϻrRgjΣ�lZ�?��ș��_���;��"qU5�M
uT���R�Sa,��5�~�@��2�|(� l����mu�q�7v� �;�����ͭ����[S��<�X�� ����W����ԃ�w_:

�CX��?���H�qO~���5��Q��ס����"�]�ҵN�6C�\h��or���Z���������gs\�+Q�Wr(�c�]u��uP�C�P>��F�D c�)���$H�EyD;?�b����7d��3��_c'��qEqO�E�p��Z6R�晿`���M��%�a굍E�u��#i-y��o��&א�/_�\�U���Ʒ�?d��9(Q$��0�\�j|�]�<��z5e�6L��ݔ���%�o��:�?c���Vc:��G�����������b5.�uH���h�)H�۔� �[��~��&0lxۍ��9�s�Y)(�|Z�m?��Y���W��[�y-�gY�b��7�$�@	uٜ���C���\N����ڰ��������c��I�fsJ��&*�f������%

��0��5Mhb�zl:{��My��!744��J�z�*��j8�؟�Ȝ�����nX:ķ���c46Io�n"��ۅT�J)O��򣐴����Vw	�0G�Y�u�b�0��O��ƨ[q5�n�Е}>"�톮L��/��ߍv�y�"�C�Ǽ�h���UݻP��W�oY�T�5�s{��P��%�lx&ph�7{rZt ��w�O��r�)o�j���7c�&Oc��)"�+�����6���.�VF��nS�j�u���ق�,�I��=D�&����֭���f)�-v�� V	��o��̲�z�m�P�w
��L�����YgqbW�ƻ��o�P��y�o4��r[�H�@9#�ѹ���\|Sw��� �.�(v4,�LSY���7ɔ
ұo�y����Z0��/�jK��i�x͂�S_7>$1P���9~被R����Ee~�Cf#ɽW���ӓ%b�S3��v��CX@]C_�Ŏo�֧������� k5WV!���u���BʇX�җ��Z?�3�z��7���fJ���@�v��Y[�F]1W] ��Y�
�*�����_e��w����'��=-VtbH~� Nռ�GhZ�􈚓cFJl�$>Q����@�s>?	oZ����i�<��;�^Գ�69�v��Q��孝��^l�PQ��8���>H~�ɚ���kG݇��MM=#V6g�`������05���⢍�9@,X���̒���Xu����`�<�$�f<����nR��n͊F
��IӅ��w�??T5�UX�KN{�+�g:ay	�Tշ�WD�1Ī�r��Cl��仧d]N�]gz,�|P���?<��w���8�~�h��?��9��Ñ7P
���f�+7�~�|�F*�����E��E�
� ��#�}�O+ں7cz�J|���0�i�n�-�~����t���eN���v2 u��N��d�-4��@nN�%��=.�pq��w~�Ҭ��)V��;Ӵ�:�Q�%,���J��硲�ؑC�3'�{�0z��l3�EUA��@�ʥ�!�h<l"���B�Ł��6~K۽�ۨ�@hh��)-�I���k]�(��A�q���M!(И�؃?�>YI֊jR�R���<޶����/���@��Ǵ[���G���i��M�#��J�E��o_L
f0�:Խ�<�B�׉��
H�)��T۝�*l�f(�V�f�q���JO�?���hĀͬd�ćXnV��e�/��{|���}�Nzw�$j��u=e�M��r\��k&H���Ѭ�n�p�s~�Fg&��N���٥��ɐ�7��6�N=$�f�?��<F7��V��zF��Qw�#���s^6�D�>��3}]�zl$/�������xwwx��50pۨ�|��_�������v*8� ���8��!#��V`b�iHB�߈�����6EE}G2(�U����_ļ����$9Y^�zbª����g�?��y�2�ݗ�[��. v������AQ>h�⦽����v�c�yo?������ߛ����z�]��)n��+lI5�K��:RB�5�z����|�F���5`m����EG������9|�aeJ |V<p�� �O��Ի�����l��#�!5����2������u�Ir���\Iq��W�Y=��1��HJvD�fC�l�ن��^�#̍����g��l�:V$����<~�s�_�E����^b���Ȧ�G,�	�ܐ��@���w���~�6m�3��{��A1d�K�Rk�^�C���\Ͻ�9��j��y�]�k�Z�`d�nd��(oKIT�IIW��?CV��k�ǫ���cnT�����}�:�8��H�%eq��C�b��(��A�`��V�����8h�vڭ��F�貜����7�bi���up����H� z���oUz!泮f�l2�"��B.q�`H��F����6�6y�W�� �w�*�_w����3�\��T�	����i���O���"����kJ��]�ѳ&6RA�H�[-9�������i���u�����j��u����>�Gm܊����	2T��=M`���`}Z�������W��HX04Վ�y=���pv�-|F-�L��[��fYw�Wx���������J2	�d��� �?��������\�)�O*C�)>�^u��e�PL|Sj7��q��Wz�øOe�է0Jٍ�8�9oiE�oNrw��z�'���dk����/zݽ��7H����zZomt0wxx	�b���M���³�Kui��UMߛ�B�\:�o$���N�e;�h����Z��Z�N=��r�r���-��'&+��$*�F�C�3X��3"�ӏ(�8G�*���c.{RV�/Ζ�L�2c#�=E[#�\��3�	�8+���Xu���v���0z��Ss�n�!<��q�o��e�kg/��$��5���L!�DUW��IR�G+�T��`M}��?����Y�ul�T4K�󪗬��ʐy��@�RU�w��½�%��5m�5/�j�:4��ģ��r�F�5��n�f���OC�i:~��Z�;����  u�]	����xFC��챶a����$Gٗz�~VnP�J^�KEHU��u�- ��sR����2?�b�u�8=����䣍t����U�׬�=�"l�Zʂ{24x��/;-Z"��1��r�u>���P��a�:9f�����.{q�ވ�t�H�f�ݮo<����X{K~O�/�T���w�yx=]8q�lFզ�`"sX-���ڽ�M��l�z�~�5*�q(�:��uf������Fu9��V���HRإ�p@�ؙ6T�Y��Z�G)td�?�HRh(�F"d#n����MQ��L���o���;�vF�
�����)zw#���+K7���G�K�
��t���kT�z�+�i�ɋ/�W5�
敍�@��zss>.�(����*��~�BR��Y
|ёظ����+����M�w^\�ƺ��V���O��K�p;8|������v���`T�ha�7{�юBI_WO��pu.�J�R}2?��|�����4�^��\y�?g !e�J	Fz鱨N���(�s��oë5G�����'c�wʙµ��+#���w�;w�px����̶�����?'�Mˏ���o�y�jT�J�zE
����}#`�
F<�I7����OQ��.n�'�+!����z �7Ul��1�?؍W�[���ߴ���:�~T����N�bߕ��"	�����Û�Ŝ���Ox�Fs�Z�WlȆ�,�h����U1�����b�M��}RCv���t��P�欖5�©�܊΍j��9�lO���]q���`���` �o��9������3�Pmt/ NC�?Ê�cr;�}Ch���e�j�N1=%w�&V8� ��s]H!��4�(ňv�z]���w��P�V��;%���was,���r���(E�"A����\zݥ*ּl��T�ȁ���^�dmlc��ǳǦ�L�nc�rY��Q���@��;r�^<FF�hD�&�Dsގ��CKl��W��w�<-��W��|�ܺZ �+�3�4�{�uκ��G�/�v�-\��5�|��CN���3�^�}/ѧ�������H�?T0�?�loJ���'��l��I�.����󲊰h܅���iV���w3�*U����¯O��MF�>�J�y,{���d�I@�x�Iab��s��oa�T.sX�zI��&V�R��e�>k0?�`*��p<q�����
Q��8�4�Zi8=�Z�J�����qV^VQh��-���pw�k��Z��;���\��{�z��g['���3G�)%���Bo>��=aZ�Y��D��)�J���̵�����K=;�g�]0P@�?3cG�֏��%"w5گ�����#��J�Lԑ��Q"$���^c�Fh*����v�@6����|]r����=O�to����!c�����/R�R�%ςH�$�Īn�9��'4B6t�TP�t��piz�FWfj� Γ�T-P�4xRN�)0%f�����,-Z����&���|��h8�h��Qg��i�4��9���#�����kb�(|`���#��g>�Cu�J[�I�
����@0��-���@��o�
��Q������WC�ťO�{R��)�ˀ& !�	�B�U�6J{�ȪTt�Wualފʈ:@:�)� ����z[//g����M�.Y�w-w��_�&��}�'��c?QWZ�uy�������~lyO�'�õ�EY��fD�S�C������;}�H!X�߀7�3'����c��ϗT�\_܀� (�mD̏6�|�A譬���j��� �3�>��6wD�,���t�7����FPU)h�|kҧ��o	��9�hq�w�?B�[XB�_<ƌ8���?cӲD���<o�`ֆ�"Z�Z�}:z�vGmH���S���m_N����;�E��U��CS�����.�Z��#T��y�@�v-vP1yv�5�g���Y��x�us�2�U#c�ܝ���]���0H��F}�Gz_%����^��I�8�"�㓿Q�7�3��Y1���R~�����3��sج�I��:�HaoEz��4"K0�)@�2&��2d	X�Q�K4����Awg�0*^v"�3����p�:���ޣ3�)���/��j/W�*T�&�{oQqs�Ƀ�p��#?�d9GK�^��k�A����b_A����ҟ�RHP��N���)��_�,�Y����I��O�[�tÑN�;�9mU�w.X�´1����G@_8�>�o�����/�}���pGwg���tXS6��X[�!�c@��P��=�� �����f����bA�&s�@t�]���w���ƣ#�e��upE�ĳ�r�PkVߜ4U�{3���T�E��?�Ir�����6$<�Y��6�w��A�d��W��?���;�����G��HX%r>�P��첷�g-�I��y��9~%Z���ڔ�
E�%�Q6>B�#�y���պUx%w�"o�Ad֫�>NAh��i:������PF��J{�$.J�מ�%�'��S�񩯯��8m�i�~j^�s溟�O��� �Ӭ�oM
(=�������sp��L>n\�1u�dy�+�W����L1�h�1Q)B�X,�I�u��G�9��,C��UI��D��I���$� M�.wy��O��}]�|BHnY��+�ӐN����)�(:��FY$�L���I%�I��PG�N��:������G\�k��������,>����J�,�7��v���62�t�%9X9���5_ņo	� �P�O��M���,�_]�z鱷KJ�	B��"^��}����,/�DN�{]�t3��_B��No��	p�Q�/.%��u�߮��30���F�ڛ���D��I����"�0�Kitәp}@'T��B�EIx���qS���^�F�iL��[ѕ��!A3ǌߍ@-��
�(b\�RZ:,2�Y���Y:�W�7�MQ�LV�v1[e���6D��K�aXS����$U��*�A��('�g�E}C���4��l7�����v�g��G�0?b�匞27�&0\�'p{-��CrG���>����@�u�=N��.��ajP���� D�N4Z�g�ihD��FYQ-�u�,b��� ��Tg+}����[���V��ǯ��cO��m��^����w�T)9J?\�0��c�`[��2<�$A���G�"rr�$�ӳ�ɑ���jk)k���ϴ%�U/� (	GL�$�t5��_ۈ0����0
�����S����켨�O^W��Ŕ���7���׆n {�}�.y��uc�gV�*�A԰��_Z���c��ڣ��20 '��TA<�g����f��&M=��XF�q7�������C2W�`����!�nu |bw�B�uz>+���`Ǻv3_����1?�'�o�Oʂt���i�eh��^�i�)����D��	��q����(e��o�4�Dû����ʌ�W����Ns�a6Y��4�l��C�����Z����S��6A�#Q:�\���0g����X,�m>�2�34��'Л,�����%��Ζ�׫�P�i�Z�]����W��X,�70��I��)��r=�����=\W,����t��=�z�]+�%4�����V�N��g���x� W��*��a��S?��4�;�d��m��jP}�>X�����&�U��C�pJ�`'h��t����r���?��i�0*��hе9
�'��qk�ɥ�؝��P�4����CZ1D�i�q��<�RRT�����UR����c�@HA�d�ɞ!�g�iA�bc�o�h{���H�O��x(����3�y~]I�h�O*胉��m��G�Қ�S!���Q>y��ȧ���A���c]�U���W>.�_��|��A� �*0_|1!�ꑊ8%��)#M�r�EW�r���#���]�l�n()z���\��?*2�����ؕ�;!&�ux�RI���Bo��O�a��0�����TI\���ҽ=�lS�]�G����jI���%F�$7�E ���.v�bi��o1-To�n0�]!�EL5K�F�׬-ߜ.5�#e?mWFw�?���-��
tHK���aa�9��E���mZ�E+<�;g#�w��w���o��zKz�HF�i#�h� ז}U�9sK��X�(��P$>2�x6D��f� S�S��Ӎt��-g��`.�,�
����o_���v��G�ՖO�����u����� �1۫����������@F�ĳⲯ]T����0X���F��J�)�?�$�:�{o�b5f��+�֑~�6����W����ҧG/���*։������=�2Uh�W�3�&�JW�����Po��;-�Bwb1T������x��+� �樤�u��}=�^�F�MH��I�����a�M/����%��%}b*��ޟz({ ^)fo6;��8)L���*[�tG�y����x ��$!��Cy�.f!�W]U���+t������v	2�����5G'�8O���&)Rǯ�W�I�w�n�gWɯ��"/`ӄ�+R�PS��e$<��7�K?/�p	f������jҪ��P�EE�ل��A��5���VMeҖ��z��IJ��$�9�{H�����ޯX!��9ޘ�y�n���;2(Q���%����L���oNeu(ۙ��z�輵���h���I+��_�k�S�>L]|���G�'}L�~Zn��֨��5�A��9{ڻ�!���o#n:9��|�������Œ��<�}��"����zi�Y��Q'i����<�I'�.D����i�X�
FFA������q����T8Z�������3��{�;��iS��^��-���T�m�LAC�x�F /*��� ��!G�>��ҽ��q�5<BݮK��>/�B�$�?��~4֍�����Lrt����|mָr?'�o�zb���.t�T���%b�4���y}c����ҝ����s�p^>6h�M_h3��D'��Q��!���w�,�e�k&�q7�C�_)/�4ou�l����j�&�1H��}�dLL_�8U�T�Ts��g�X�%�gjἔ� �/����6V��)�z�u�A��Ŧ��u���e���|�M)�#�/�<�͊��Bi����~��^W�t����Npww������=�C �	���������ݿ=w�ouU�:�n7�4"�'Ї���뎸�k~M�em���ND��з�38h�n�v�Atx�N�,��Е�g���:����y%�=%mQ�f� �?(`�(,�����Xs�9Q������MK���=����h��緍k`������p��1�i�lZ9G��6w���=�#���-1@���7d�'�-���{K�&���N�i�1yu|�e����y҇*�%�ѻ���Y�`��lW�Y����nv�9S�yCo�3��	)g�#�U���D�L��6�w�s 84���˽/Z��5M��M�mB�|D��U?��D0��E�xp�~S�����U����9��y{UU����Pb����AAͳ�@E��ҧ�⍟��F�))i�a���q�\`���%D�q�!�V;#8����i/e<��:�m\��rQ�I	��T����[ZJ>�uL7%���M�:���S�;$(�M0gt�DU��'�~(���!��?e����0�Qoyf�3��;�u�w�~��֤(�0Oq��/��Ql�b�w�k���\9��8P3A߁Paq&h"�$Z���Ո�Y��>�[B�뿋W�Z~��S�v��Y�yb��Ó#s��`��u~�rt�\���_�JK���3F����Y��~!˓����|3*?B�Qx��y����F ݴ���)��l$dAIC\D�_����g����bq���')z�����z��E�z٦��_������%p^�����G/�P�Û�}i�u���`�o�;�����g�}*ky��t�k��yơ�MT�z������I�}��@&�k���d�wXC�˃ �O.8��ۺBU�q�l�B�J[���i#0E	�S�7;��# v��~��C_{!A~�U�-nc�3R��A�g��ΐfnp�������b��P��jvx���{
d�������A!u�/����ă �$'m��l��b>�J^/6�wo��?�?�ضI�݅�8��y.�ړw'�?N�\uV+�1U �'	k�g�<�qj��nFdO���Wz8��5�J�T����6���<���UO`��N��z<)w���`쨣����F����ŵ��g(��)�MOJ��8��)#���<���������`M(�����k�����Ӂ5�	3x
��b$��grj��޿j�ab��S�{
j�sU-�j =6��q��o��#�#�^�њġ���ߦ��6�ܑ�#�zk/'��8�3��\�@2��W�?��!��w�J�AS��B	_qas�4!�-�pr�����q!̾�a�3������ʒ��^U/���N�9� "��l(�)*�b����ڿz�U�"1�4JP[���Zv6�f�<�;wGZ^vL�-�8�~���˥�(P4���|�pK�gO��X�������7i��[��S�Ҩ�M5�M�R��ޭ���v�f4o2�/�ٔV�88`�K�;��Q7���*�d���kR�D0��5I���b%#Gowsf�Ξf��V�ʵC��U��RiRh9gy�W�r��0��~)<)�����h�J� �{�S@Mc�rr��zrȈ3;����w��ڧ�"�a�i�rX�ÿk�^+�f�� ]�qs�w�Ƅ޲�4?�#ȓ�>�=���P_�Qʹ���`$8�c�,��7L�.CJQ� O�qԎ��m8�zm5B�<O �7y�Y([�
��#nKg��o��+��$0���ꛆ`i���D-$������w7��/^�PgG�9e,�y�;���˪�@����ٕ9�p��K*w��9(��Cٜ���Z�h�I�ʝUoJ9=9$��Z'��F�Y�@��A�y��]�x��V�e�}�Ub� ��^z��د^�� �k�C��8���6�����;���gV��k���M�?i/�] �	]z*c�5�v1ûdT�S������Ru�I��,�e��3b\R�����U�5�"�Y'B������=��him�ϓUޓ�7.���� ��Od~��,��'��.�5˼4���y�y�5��O�~� l�0�	Ԣq��JA=t���L6�3&!�ŗ̆YpSD��g"���(]O��������[�����f��S���0_Iڹ)�p�&�*�u!�wny�ԯ��}/�dp�|T��?�#G�d.��Ȼ��5Þ�ho�i�j|0̑��G�8Đ��РA�Nv=�[&��#��)����X����K"��o�(Ef��Qd�&�m�ܕٟ�����@$p����&AoO�}�:��3r	�7��!B
���d�؅���7�\���gB&�=7�E>�K�/����ģ��}��#m����`�o�o�����ԙ��F�FB���$����K�$�Õ��c{.<ۚ�q��� �E���GZ�8}�Cǥ��ۏK��H�.[���o��&>�6S��X��n�O�F����M(����*������p��� �z���D��弍7^D(I�1�����:��L�Gz�p��<o �0�"��l��2t=�2��俿[��0�2��`� �|v!X�CIfB��2��F�or���S� 瀃���(��Eȶ�Z9��I�r��%-6�	���'�"s�a�|,�� n�B|����ޕG��`ԁiU���1��?�%{��r��zs�X:(&�����.5�O�E�F-��Ik�p艈*b��a�B�+�<N��N�sχE$��}-t��<��I�U�C����3-�/8��	��-��aG���2[����kn�1dkF��\�� �_H2
�6��b �s��,��:D�
c���Z}�\����e_����T��:u�}u���I����_�:?��R)�N�>�9�qxL��4J���Ki[.�'jˇ�^��k
�ϻ*ŕ�M�ۆ�E�d4��ǿƨ�<��<��$�J>>�*|"��ۃi�'��R���I%"4�Ǚ��:�O�Ț�u9Z�}&z��ʢ�� rv���	���ڣ~����/@���1����Y��'�ޱ��R_��un-ر]�hXk�M���y ���� -r���8��B��F�������US�T��wŘ���C���u��"5��m拞�1���b���.��jk���5���C�P)�`n[�.��sުl�7���~ֈ��izqa��4�oձt�.k(�o�/�1��5D��fn�^;p�A���^<Z;���N�X���ܚ7{�����_�����L�-5|�g�h������6��9�\^��yo���N��I��<7�;zKN�b��oc���E�D�Fa���!є��w��Q�A��P�)��Z�͏vD-��k!�/�9���!��h����H���-I�Nc	W�@����WŜb��8����o����j��>�^":� �W΢9H����i�B����R��W�g�#� ��$"4�#�c��o`�EE$�j�;J4E��Ў���BC7_J��|�62��X�=<<�<������;\<U;��o��o�b�P�	l�3k����rˑ�g�����@�d��~R)I���絿zm�ݕ�*��ܑ�ﺖ�YGo/��FH7C������ެӓ��Sw�>n�q�*�/�b�����ּ��E��h�An(�N޶Z��_���v�u`c�PlG%�z]Ւ���\�/oW3nˣ�����^�tnxY�e����M��-�o����ᑽOW�
��)�6A�_�������m5{K�c����AG���l~\��;��
rA�	O�U�LۓL�+�Z�d��9-�#��jµ���Un�3]��H2��|��<v��P��Vb�ה�͋��b�#�cѺB�ˢF�	�ab���{�c0Mǌ��Qgfv�<T�)/casuvB[��;`��{�~<��֒|��?l2��2�m��@��^ya�%�FB�a���M`|�ԓ��5L�����~��@^��t�<�ǖ�*���h�A7>����w?R��kxz��DИ��QMS�_�G��%{��-c�R�󎈲�p�ȈO/�a��3��s��cky.��7�G�b#�r�!��	�nxW�)~�y��s@��1G�c��oӘ)��`o{���s%=�(�o�,�x�7ׇ�i=�z[]� ��:�&򐹂���B�˼�]�!s{�ݥ��ݺJD����i����:a�����,E��ߔ9�;jŃ�} �"�xq�q׎��J��fh�ޜM��e����M)��hՎ�����ഐ��M6x���\�.	��S�gh�A@.pτ�9���G��A&�?��	�A
X���Q!=pz�7-����<���k��A�pK\��m���6�rPt^�s����q��k���V�7�]����I�ͦ���l���qS*��� ����T�
�Ɛ��d!�d|(�sz��k:U�qZn�Pg��e�'�dgf�^� kN:c��`��<����6nݐK��8�����n��To:��=$z5��A�}ga�k� 6D.k�*����Yf�������ެ�&�ފ����m�EWc��"�gb�H�{����-�O�]��@JS�-�oE�KT˺10�21��w?�N�#�[z2�J�9��Hwa߱H��[�a"���<�����w�:-���G�t��}��4�_�g�`7�J��X���$s�I0���1|%�5�
Q_=��RH�^�c{�y�q�:N9`����ޙ�ž��gw�Ȓ��j��>��"����I6��uE��ͬ�G��\(#� 5�3��P�o��uLǏM�(�(+�����&���(Z�LS��'ˀ�����*��Pa!o����esF@�KY�&z�����;���I[��*�vx"@V)�:� �a>�Js������޷��\�1�C���tG��!Tc
����So!�j_օX�Թ^����˥�/.�b�O�N��Am���v�f���r ��,����TK�dp!�f�j�nD1�lt��5�1��^T}�:} y���l�M���f_C��С^��q~�
�{�q�K�֖���`?����`q�j~q�j��/���^b�;H#a�����%�9�Y]��1��nSn�UJ�����X4P�Gq�ZZ��ya�m�^O�ӯ?Lb�,��0,;!f��ڠ�s(&bt�a���of�7o�v��*����A��t�D�V3��Ȃ����W���u�}tp�g4��Z*�G�(\��i�Bj7sF��w�(2�>}<�l*��̳p�����3��d����k+�P��mfV�p3��e!��Zu���"���������3��K�)�c�X�bNI��R��H6/	�(en#��� �w���|Vc����?f ���0[�T��I��t�����9�,������E��&�n�ޞ�G�;�E�w�A��5��;�����V.��=2��`]�6Z3�kl4 �ba�v�|�p|=�*�G�/xY#���t�"�u�i,�~��n����[k*Z�ps�pQ:}rȹ/����!�8� V��錍x��e���PLl�9�۳��}�@��	E�����������\R��/#�OL4����m��ȷ����"��DJsD9X�r�-�{&����5=t���́9w�����\L[:.J�����,c�X �و����Ȅ}��h둭��=�Ɂ^v���x��)S�+ܶ#[�Ї)1���;V����}��;�%Hd� ��m[f���5>���=��Jݟ�ǳ~��!
.���1���f����R#ok��V����D��s��6tP��1�+�}��Y	��_%�;��6�	�-��a<���>H��+vX�M0F�?��|? Q��./\���у�	5dG%`.l��K��=���C;'��N��y�]̞��Z!/�3�W���-�y3�~`p�x��>xn�<��n�J��9�"��/}����T�h�T�ς'�����}��Z�7'2g4[ȡ��ٍ��a}����؟~9>;�i	���L��!�G�Ϻp�����@�� 뉒s��az�'�_Y��"���k�I�a$;��;�7@fj�������3��:턜/�ivo������\������w�a2R'a�u����oljbCh55�&$��g��V���b3�%4����s��H���A����6W��>E�C�ݙ��
���2G�;��-j�Juɹ�@����ɧ�Y(>uCɟ��xl��R�Z�LQ��Ћ�XNC��m��Z��gʐ��mu��a�kN����^��S<й���i��k���bRTK�8c�󘨎5���G��a`������uo�+-�ٽi\ؔ�2��bZS�<���ZJEi�D%�V6��t���itҪ����y!8���7W�vynm0+6Ǝ�0v�|��@�8����&J����]1���i
A�+4uA�,/��x&s�$s�Y�
�}JZS�}	��z�b�nt��şA�����R!ǥ�U�F�o:sS�HbFn����@�� g"1����Dm
���1�9��m_|t.���Ц߄�����i}�ͭ��I���_P���8�$�x :6�;�4��e����-�/dk��+�i0��E�;%��|JN�+��?��;��(b����'"Z���%	s��.@��LBY�*�zk���<��~wj�v�0�''4-�h�{���F��(��f}t³〵���ʽ4<S������#b��_o
%�x��Pd���r ��%}�^,?��$� �ͽ���=��P#��P�%�:#r
�3�Ey���C^�">��)�-Ti{��G=�S�z)љ�+��5��~h�9D�#��f��$UMq=.S� ��Rg	����Q��^eM������it�0�[�sXkH��#KT��� ˬ��"�z���2���S�Ի_�CYI�N�2N]�D����k��k��2jt�̥�5���}=vךK��o��I��D �v�����!G�I˝k��
�>�$qv:�@��B��� ��d� ��J�֯�ž��u����&�3�N�1_3�?�V�L�;���ة�h�E�? Iy/6)s�(��6)<��hW�0��b��~Y��X,�lEs��Q�נ��!.��CK��u�Ou�������h��ć�"�'t,����˒X�s\��L���	��}�n����u?�ϳ�G��9M<�W2b�Is�OtK��f�M��<�x�Vg�ٳac��~f�7�r�l=�t,��ij�̖_6�Z�b`�O͹��hx��7p�	W�5�x�����c������|�7-�����nś�(�E�Y�>�4u����������{nT�ĕM��}���}�6�Ņ���U��P$���@Ev�O`����N�?w�ˢ�i�Q#ͮ�3�]#��K�R�C�c�o�D�]�͜��#�ß�Yc�곐���77q �����>��R����۶��Ɇ�C�b5����6|�	O�����#ս��5m�>�����e�O�(����g`�;(��|�Z̼�هw_��|/����%�ú�o`aG��v��S�S�`ݔC//okRn��kf���ض�J�/��J�Y�mi���һ�!Xw}]��u�y(�L��mk7�S	;�����r��.�l��%��(e@
]�j7m��6I���j��4c��#.�`:�-��2!(�$�6����}Ӷ���Q�@x f;�s[���^p Yo�@ �u�Ї�8�y;d�|��3��Vjk�>����̄L�����r>7�0�ڃ[0r�-�z3 #�=i�k�i����0����Q�������N�|`���B̱yĻ�/`��f|�3�*2����c�4g�@��V�
5�v�t��{ow[~t�Y͹�ԦC1��<|�ڹ�^Ț� � ��Y���Ԝ=�U��:)%4Nְ�\�I[���*��Bff�7�ٌ�>�@6(�L����Ԟ��i��jN����]|Q�ة��e�?�	%2��}x����0lNk�۱c�*gn��}�a�J7�oy�}h�.��<��y|����r�{��dY�-_�u�L�!�e�e�<�=��y�lT�{����;�ỽ�e�I ���%9��{���c�o��P���Ù�ηm�D4r��^O��^~���s��]��3�d�cN'-��#a�	�<�`q�k[�[}�SCpq�yȭ�VK8����Ý"��[ͼ(����+La@���^���!#*�C
�"�,C���[�����O�^����ˆ�Y���H�ͽ�D���H�iH��4G ����^l7�����s7�F�N�2MĽ<8ź��i��k����Vu��g�f�k����L��{���AV5$V��ET�o*m�q;�����[�o���?I|��B��z�̲������[�$�n!����� ���g�
������)z���pSA��ğ��a��k����X�3ߐػ7���Jd��6�fJ?�F���Ҿ�#)t5��y���(����ޓb��r���^�1�i���_l:Y6�1�h����*�5k���N/�N�7�"I�=��K8p�L{�s�@��c��j���`�\�Z�;{i���z�zU���%�2匯���wyn��t�q����5O8���Ek�i.A��:k��@�o��Ε����C�|`�%j�,��%�"bQI����ǉ�}i�ӹh�*�Ǚ�%�2G(�ON��K��яb pض-��~w4R��L��t�Bn�z�H�v-���h��2�����n�j�3N
�Z@紱Oo��p�~���_��*J��૫�l���_X��%b��A�۾�_D�;���U�Pj�/�l�Qh�i��j����Of>i�bd��i/EgԶ����Q�X�9 �-���.��!/έ��κ�v �vƠt�x�<{ ��?�R��b�D��XPu%�)eħ_X�5$ﯗS ��W��%���{�z�x��j'"����$��{���qca�tN�}v��\j�t%�Y5
� 6�t��D��9�Wȅ( J�z&~�uĽ�D�����EuOC/�\��S��y�9������96��|�0 i`5�Z���e��]=� t*�>9���_�V�����r�4�AK=��59��%k���L`ŏ���/K�A�֒��p�'q�ہė
�\s{���z�+���jb˃6x��fC蕄gjn�+Ľ�N�eI4���+3�x�5���_�6A�,W�a\ne�!����n�ژ��>B_�?�eW������O�Si_�R���R���r�����3�kh��-Ƕ��/č�6'G�R���M�TH�D�s�Ӌϳ*cο?�-�X^�F��,��C�2�$] o�^2����#l3�Q�t�Z^���\��R�kAK�̈�(l�vD1�x��"�/�F�G��p�C��dCwC�3�\B���I�N0z�k��b�`R�Ͻ�s@YI\�-��:�J�Q���Rј�2m0�0��֙�-���h���F)�� Ϸmɏs�t��M��E�1�_�̺�"4�Q���(�����T��#�KO2��t*ٛzAQ�Z��^�U��"�02�)�����]k���N���ÎES`�wk�,�6X�-��
�����Of�����Ūf���=�ȡ�Ccߤ�Mn'Y"�n��ʢ�M~��q����%w�zG��%j�B���6Q��q�s^�-<����&5-���ߩ�H�bq�I�_������&�������. ���ձ)�UpC;��m���N��C8�Z�m؞�B����d� �q��}� ���E�����!,�Rw@�"�w�`�c�� @��A��<�8G��L�q�B��'ą!	�)[ЧL���_\��=�z��٦���j݃ڔ7J#��_�g���&&�O~�|����9�m�BlZ�[;/m�8�^�]����;'b�8�񶘇h�l��_�1ѕI'���a��M@�F�C�w�39[]�8��~�Ez��Y99kG[�v=F����f;�9���V������������ ~pUW˩�+�����鉽E����WR��a?�J�r� ��s$�;���C	�60��ڿ�بn��� �c`����ԯ��VVVQ��"xƭ��0w|�~�4��np�(�֪��m�o���<��h0Dv�N��둂f����o�ou���!�w�� JJ�*>�5�
������eP��"�0�593zt4rI����ܺr����=���js
2�ۈ.�Q�"��������Z�S.����M8_����@C/R(���'1>�#�mn�G���᠕��������	/�w��_w�Z<��������w,����A�VPP��;�l�[KKd!��Y�ОT_����*-++�fΚ�4���tǍW� �uv�ȥe������FةΘ-Wp���6���R�#K�B�������ڕ���	.�l����A�O�	;�Z����ՙ 0<��4��;8#�Įc���u�P�$g��j|<�4?{�iD;�dQ��w9 �z�g��sI�>9�f���]ėҺG��#(]X�}��O��Mς3�?�0m��~i:��$�r�&���E��d�p�U��4W#�(<8��+��
I(��J'��s_)�淤�+��(}܂�����z�y[d
N�o�6������x�ÒȄ���%�]��j�?3Z9�lbE�٣���~����[��-�ȥ�����w�e	���!��tU} ��Q�'��B� Z���6�Ȏ���=��xdp�w/��|�A����L�<��s;|�8�db�k�j��l�tե}�Q	���i�*4s;��S�0�ۊ�xzhw�ܳ��$M4]/$Ĝ�'/�����KD*���y)����lS��I�p��˻�"*�:� ��7�~>- �!"&��C��0�:>";h.��V��tN�^�-���f�w��PB9��tVEO�Xý��L�U��"���R�7uJf�V�AꐺN�*�MO��s��q�m1�IDS�&�sR�L���I�I*�0l@�=5��:��)x��P��y�h{�^��{Σ=C�7��[꬜4�<�5uÈ(X��]#��ªΙ���2�.���r�N#��R&?>a�g�#������k�����U2KT2\"�)�
;?���, ܃)�j��)A���>��M����:2��-���B�2.oS��')[U����,; ���L�4�$���Oy�)�R
�4�:W@s�n��0��\����������K5\.�a��+�7���#,��&��ҙ�2�Y^�
fs� �.~��-���P\�3�p�#��i��c�W7��(�����ԓМw˷X��C�\c�'��h>�E��Ov��%x��X�5�0�m�=�)φ��K�7�LDPS�&���H�jul,h�N�إk��j��\z3K��<�oG9��4xy٭�j�4�_'��=[ ���؈�{+x���cЉ_�����2d�z��ni��z�����o}��J�����#N��r?���xx�	Ia�|�wmǅ �גQ�
��;��,�9/��Yt��z��Ź!�d��ъ�8x�M�/�+������S�������I���uq�4�-�!}i4�j���b8�Z�»�׊覙���&Z�
]�`R�$��9�|�S�L��4Tuu��>.e��~����>3��}���ʑ�s ,��qH�q��4?z�k݉���:��~5���!�3mTc�l�{9��G�����/�2i|�E�[��d&������BJ7��l�#�	;k�D�g4<_wH8$,^�:�$Xgp�~��L�|��@���3�'�5�1��ٌ�O�G�9lm���SӤ���8�~�K��4E���|m�9��>�����ћ��)SuQ�h�񰏳m�<_���Z�oS�s��;9�xr�U)�ɜ��4�3qv��^��2>S�g:�G�r��O*Q�K���aZ�^>bpMM`���=Av����0	����bgŦ��máÂ�3J�2�12ǦΧ>���p�:̗u]a�c]Ű���z�g��Tš�U�7rȰ(Q2�/�f!��p������E����!N��/}H��(�oպ�
Ʌ%��Prf��W!�:	�`@�Q���OMp�#✂k���~b�@,�n@���5�V��z�>��TV��q�A��g�8:M텘�oHIy栵���
��Y��mL��R6)ˀ ����{~�r>r"�����5�&�h��͑��T�Uƙr<�׷d�ҽ��M�K���u6�}��`�Ju7i?5{��TO�b9�9X�Yw�=� �����Q*��]��	�Ȃ��n��@�I���G��xɸWNo0��G����3�$����Mp|4�%��KO��7~�˦�oy7����S4$�.�[ǎ�l�]���6Lj�r��T���i"̓�W}:�p����b���Q0L��7�L��5�7���R�0��<x�Y~A�8�2F �ɞ��:C�{�h)8�	�ݦ��9��I�}}��կ�צ�UqH�e���H�ӟB�{��	�a]LtX��o%�B��-�,��������A��$+t�#�^�1�����/D?��j�%�B��Wc�p��c�Ҟ�w!��h�Av�}���7 =�ߠ��"�C@I~j���{�-���5��f��LC����hȠ�Z*�����$��-�j���5�=����*�11�ߗ��9WW׬��%�T�����>�iw���c�vtv"���.��u;��ܽ�Oq!���H� �T��}�f{p3�;���;/���G�z���*c�ό^���Y�࡭�q� Y0�6�N�����lgA����=4��l���'r�m�	�J�N�i_��\�A�%�a���#�Ll�e)��m@>D����W����^�ty���g7�,.j�'!�����v �o�� �*��a$�������_L�3Ng����i\�I}�@03���Og���h���$,$���NS����v���tc����% �yt]@e?�o��[`%NV��]w�L����a�4Tm���}G�Kc� �:��zE��8AIA�X��<�a����/.���H�ϣkQ8vsQ"��[��O��!�_=�*[�7���o���6��r�?/���L�hB̙[e��F"��-\�F�#`F���j?l�;�t+�T��|�6X�n�8�P��}jUנ���$G}���*�Rm�>E�W�n���>Y34ĵ�=��/�g���r4%�a�b)	�@h���K<������!���N��8��P�O����wOUS���<����l�,=��5���e�c���OD�������յR�t�J��l�㮬lT:ޅ<J���	�ݜa/xyV���6�Ǯ�_��Z���ǅ���P�읰%\o�IG���������qM,�^S��ن�'��T�/��k����įG7Ď��������� ���7�u�]~�>�0GI��<���g����r���TZ�t(ߛ��;�e�g4� W�0�;����㥸�x
�}���%�.{,��"���%Rذ�C�2Y�Lg��i��/u���"��&��İ(��CZy��a�Bst���s 4�$G��;�wT|f�\FM�Kq���*�;6�b-��~���j}[ɤ���9Xd���F��^��W���3���'L|��
��V��"R_�%͙����\FԖ(�F�xۊ\�_����K���p�kmL<�x|~�����Li��~¿�LWÎpv�>�H��ŵx~1���k'؉iՍ�~K��c���X��).6ń�>F9Й��E�WހM�۩�H~��=�m�(
�F�-���!���5���# ��l���
�Zw}�j��:iE+R�%�f2U7�s�V�w��ON;�ZK�p�%�	7"тQ)��':��
C� X�Ń��m��2G�:?�s��_�yiJBJ��q���j��
�~W�_��VK~D�G�=�D����!�2V����v�h��y��T�S��z�� �	~àR��D�� ��4��'t�����ZyzB9ꛤ��FPK�c�n��r7+L�����s�)t��%��\�K,Uۇz���)�s_�Vp@���%�:����
N7��+W�%�s$��}��U�K~�� ���Y�뾅]�IH����8G�V#oz���ҩ~��2� ������U�{B�9��	+�b�4�ƿ[�t�wo��贼hlD?>�T�'~S�%�?�ƫ���O,����ka�ծ|w���0�:�����X	
����<��] ,D�����oZ���8���"�|r�XC�~[(k;��'�9��}(ɩ�6��%ve
0���U ���2��~G��3�JN�_�1�a<��xK����ܜ��%_Mb{�J�	�W%��'D�W8�B�7�">�Z
}\d\p9�'��u�z�Z�9@��?�f���/D�$j�p*��y:����6�*3�_`Ҿ^8mUy[˜]D���f����֖�x��14�BV'��U����W�<x��d	��^>12 ��|�h���o�q8xK�8p�cO%ƶ�K\��$1)MV����U^�d��KRG�i�ρS��k�m�l�� ���`6��im��rH�~.%�މ�cݎ�4D����זӼ�&�Ѝ0�ulq��W��%��N�eT>?q���N2�I �x�
ՑiU��Vitfeq�SEF�>8�É0 �8���kq�7��_�N~陝�h�'a��~quH��r����oM��2¥���6�޶xLX��S�������W�L街�)�ܲ9��?�M&"[��R/iVs,:� ?*�*{����f�:?�n\���Ӛ��]3Y~�d�-6r���XY�oO'���EQ��z�������������lP�(��oy�d�s�O=�*(*foF�W��1Faں��<�I�٭k:���\��` �i�cY��F2�W�������nv9�ʛ�#��~g5����)��[!c�i���-�@�g�'ާ �>��MжU[�N��53�tX�02��ޣml���1l�>�0��'�A����|�%m��;c�e�e=��9�c�&<�/�����+X���p��w����u�$�?{�}N�Jd�g�?<�[���\�2���~����S���產U!�|;2��W�s�D6��/�Cv�j��n<�KN����q�g�ծN��8�0�Ⱥ˦��6&��S@�a#��;[�,ҵr��4��t��4�x����+���>�k!�ބ�:Ā���3���2)V�yJ�9��L+&�)�WXS����(��Aa�L�Ԁ�`x~����*����$�}�'��*�=��L!@�<��*�B�VOL�٪�N��q���`Hxq����xٗ����58�w2��/%��T4�p��ʸ1��f� |BA��X�d���.�q#���r��W��Ix�W�`<#l�;�ڢ�������@�g��_TW	�UA�8���o�Ĵ�,������s ==e�_m�㱂A�$��	���vr1V�� ك��1�����y)�kx��Hu��w���c6�a�&��V$]�Z�&� G�o�a�xH��qZǗ���r�` �j쏼�� �e��oh~SEM͹*�M:��CuYd�$.d�9:��o��uv�Q���1��I���M�ޞ��Ӹ�\�׊%�I&���e����ꦢ�����1e��ʳ	�G�S��|��/S�VX�
,oU.7���6�kqz�-���q���k�n�p�¸�a���0���_(ٔ��f�U�e+��B�MT,����Z���U3�	�?FHk�m��T��3,�s��9�9�q�K�?��e�������U���Kwʭҗ�d���o�����>�]h¶�Ue:��:�mn�
s�>����|���zz�7�@�o�^��VK!��� >#w�'K
�a��M����Ÿ�͏,cTd������7S�,�K��q)u4��=As7\m,C�}��C��i�������M]�2�7�J6��ݪ�r�r���Ck;�[���q���k$���Rҿ)^�rs~�\�C	�%*�W�7;{����T�9!���Wl�+8�Sw�����=;<����H��c`�ꏵ��଎icήyY7 g�C]q�|!zݬl�h,'z0Z-��Ij�V�V�_�Iq��Eu�j��2劒�Ԛ�u�-�OAl����h�x�TY���*b�F衹o-���>��S�D�yY;��f�9�$��ΈW�<��K��_kS�l3�]Ɍܫ��i"s�1�Z�'�mml��S��B?���fZ�Q�e����������V�����5��CTf
��h$-�GS{�W]���,��A�>s�d�Id�_eg��q�Ą�8���EY��(�uJ��W�~�?G@�Cď�u�,F�_�AC�r	�9n:��_4�ً��X�l(�3�y(�wOK�4�*)�2o�)oW�E�\\4�����]��Ӹk�qw	�ڸwwwn�|y�����9w��9�����V�Ꞁ�\_��� �%V��ң�t�J�� �a��s��
ԓ�̯�+~�L�5�4e?�P���	��5LMt(z���� Sy����"���k;�J=92Cy~���D��F� kji��[ԗG�rJ�?�V�T0O��Sǒ�1j{P;���:M��E�~SU�Ԍ���E���$7]l�S����k�<�U�$yk���lm����\
wI,�r-�[/Us.OJ±c
;�[)Z�N!��.\Ժ�
?l����|V��y`A6��q��Za3S�"���.ul!r�QZ�oX O��A���X2�)�L��[�s���k�	����=�O�ޭZ��sQ#5�)E����*�B��JQ�������	M��{F^=g88�^�g_<p>Z@��DО`��o�\	�Ha�!R��N;5Y��Ұ��i��[�#��������D��������U�F�kꓜ=�56��i���;����&��a)�E��ѵ{mGE~�/(��ڷ��5�CN,-�/��jC�s�U� ~�Kʢ(~� i\u=%5�{2����b¤5��{Z(Nx��9�-_�r?{l�ϓ[���;@v�5�:U!�)6r1S64^
�ӍW�@��%L;����Dg�-f���"���^��)p�?�����V��܊MpՎ*��{eDpV���$�$fY�\�.��)����l���5��1E�����2�G�Pɓ�}Q�q�!Aݏ��򱠛�����K�摧�h3M �L�+�-ߏ��M�VAہ�j�4����|����1Òq��EU��6��**�_�����܃'�$��׺DB��d�r8��j���۽zP*���/Ѽ?ô��[�����"!!f8[���D��`��1y�\�Q�ȡ&���Ț�͙v��� Z"��[�����~�H��W |��5P�w�nPezXA�t� �|�m%c��}��.���Nˊw*4�Q������<�3�����يZ��d�rҙB������/�)��9u=�0��:���۶����ʗ�fn��`+��M�����>��_�i�ђԗL6�xuZ(a��������MI�q�L�.x\7�F�]�I��h�q����k�z�Y*~B�'��������PG��g�0��N�x�Tq������d7�,����f�wy���W᱉����<��J���B_�>�32�U�M��V�w�X<��8�%���L#�T��i`�W���b#��Q�4�[�{Y>��l�Z��u�;�S\J`�*N�+�x�YG�~��7��`���[X?q0����}��i�C�P�3�8�Y/�v�>�~��"��C��:�~Y ��ul>Y6����{.3��ۢ��S��R̻ٔ$`mO����a��c�}�V��IE�������-+4�hI��=�����4�[��D�ٰ��I9ם���k
��ra��� DO�֘_ӑC����<E�����x���j'�3���I ����C×���u%*��y��"j�O���S�c�����w�Z�f}U�>�W[_�la��>+�a�p9�hs	mG�O�E�l$L���N`(}��T������Z@}q�v1q�r�QhϚ����)�d��M8����g��z�C;oJI��[��`1S�������'��Z����a��C�����Mt{Uq��S���l/�*�,�U�jlN�Y���'��g��prjy��H
w~��s�=�����1�;��y����h�..�k��8���9�LE����)��F�3�,ꮚw��e9��6N���SXI���]���d��)[8�g�3w�Ύ�/�uH:��'������������u�dՍ�]%4h���ܔ�#x���A���ʚ�Yh������]���c	�����"8�Niݼ�X*G]`��tշ��'0���g�׺�[�"z�?�ĜM�߰q求����YwK-��y�������a�(�#׏8�7c���co+A�q,����*���P(�;���+���9%�T9�L����B_����g����K��-xV4���Nt�)��B�L.�7e8���L��l�/�QN$�h/�q!I�������(d�j��(eq���v"�࣐j���@y�)��+y���Y[X�H�S��S��
��ǋ���i4�J����b����G��q�x���)��cXs�X��� g�r]��4@��D��aO��l��p{�����B�h���wx���p-�`_�M��ʼ����K�`��~�����ڜ����zi��ޮ�Z�V�*���퓳���������o�n��fP��i�)"�\�Q�i���gئ�����\=?�`t���{��I��}�WӠH�L�,#g�S��8�]A�a���?y�<��6{O	�p)( Z����e��`80	���z
ze\x���e���iw	��d6WVlۘ���h�#�Aܪ�
�R�16���rDZy����i%GJֱ���Z�ha--S�0�'v)�f�9k~�	�H�җ��1�J�������X���Gk$(4T���G��h�Lh�Q�#�f�Vj~�ʞP�c��]�-�}|���;yn�d+�j�����xv����?�8������^��� M��y���BSq��b���s�y��m�M�oz�2>R�!��Voi��"8�}&�~ f�{ ���
�Z!`ɨKBO���҇�s���>�.Hg�)�Tj�q�gq��/��f�M-��6�ۑ%Ԡ.���A��){YK����u�O����,�wƿ�DC�0n�e>�w�?��V'��=��K����y�k�G!�<���`dpZC9�-6��W��E�߹�.D#��gЌo��afU2Z6]�[�䠰ѽ�*EM�@��Nm��dT�h�O�.�z:��S�bJ����0ϑ�����*�C�o>/2t���(���F~��DW�51����&��S����|��m���]�M�.�mc��`қLE;������L~d��	�t?�ї"9
zK��*����h'XY�GB���|�)���G"dF���^�&��'������W�X��#�0�S��ܬ�.ļ���ǥ_�i���"��"�1F�R��m!!M�굡�l=����[W�w/O
�+)����]�y�.�˼!�ߙm���6bD�T�͟e��W���H�ɔ���K��$9L��E���?`q h-�`y:w��Ӷ�S/�)/J����NU�������+�Ķъ�R��X��Z��ٴ�D�~��da8zR�yS��,���V�[Ȑ�V0V7�esx�M:K�!��7�vE-��(4��F<H�]�ʉ��s�{�;��T>�C�����A���a�1�g|>���S�F'�.Z����I��g}��]/y�3j�����D�
E�\|���W:4/6��:Ưs�m�sRlj�W�����~Y��i�|�)��_Oa&Xeh��op�(_�B����(-�ar�wTV�i��H��&!�������-׷T��J��:�a�k�ˈ0��j���+��5=�Yk���4g�2OB��@vڏY�ۓ�b+��V3�,�����?o���rۥ�'8P���\-.�RF�=��0����x1q��~�;�w	���]@��e��_���H�	n�b�;3o�4��ɮ*nL���R��E@�%�+�3�#;��R���ī�[�8)�Ep̕ƘG�̳��zQ������#�v��55q���VZ��U5�?��0K��}��{��(�~|I �E�bnL��(]�;th^ \|��n�9qv��_��5)�R��:(3�2ϫơ�n8��Ԃ?4�$�ٛsq9�%�{A��J�,�ȫY*,aZ�;#�X�������*A�?����Lᯏ�%`��d�O������ XH1�(�WU�_�s�󫦑�>1E���4a�K�Q����;�#�nŹx�m���b;���V=nJ����p+�N�A(�o��5�4�����?��]���=�t/���M��i�/{r��
�3�-8x�*�&���;����f�;љ�w=�*WmO(��������Y��
��w�Ajb��j�b��3A�ظo���e޺���FA����@1k�z�Q~ƟX�KK����g��C���������,[�4B�~}�G��^��Ҫ�O�6��ן��u�ߞ�r�'T�v�6T�q���K��^�rk�[Y�k�D�x���6h�Q��|2�GLQ�{ÝH���lQ����Ma����xO���3���K��SjĻG�C�u�dθ�Gϐ���So�;"�-\�"�ea�bY����X�����-����A��&DT#m���W����W3Mb����b�n��Ge�5����,4����V���'h_R��F��J�p��,u�sN�.�0�.��S?|q��/����'y�_�A!�ڴ�̕qڈ&��	��Ch�����E���#M�sc��HNp�9��T*�бh-��_>��_n�`�F�����^Z����w_�����2)؅��{T�l҄�1�����텵�ևssR�P&±�}b~��7����nNJو����gNy�� �/TE%��;v� ��q����r?;4{����4:�g2cgP�1���E�7բs�?v���+�Y���,π��)$�P�o�KOh��z�ο�	A�<U����/)ш�7�}��$/�X�n�;r��&q�G������Y�n�Т\��I�ߧ?,o���Ф �O��+��q�<�{{f�P}ͨ^�y[�k�sm_��KW�~�pnۯ�&8u-��{z��0N$.^f�ȾƊ0�.�ju֯�3~��ʠ}����)M P@��|�G����B�q?�_��c{�^�gB4�s>�(A7���]�eQ�*b��^^�&�5A�o2q��3����3YE����M/��M?��ra�S|,8hc������Ӿ��߲%�ݢ�O����f�*���>���S�Y��p���}��B�;���Wi�(��I�-�Ґn}Eژ�e�T���f|�s�F��c�*�A��s�ALc0.{t�SF�%8�|��I����x��wիL�=��4��ͦ�W�+�9Wt[��qq����K1�S�lٝ��S��32<�ޜ.u�t��ٹ����&4Ҍ�S�R7����OUaˢs{�1����7�u%:�����ъNGN�������U{5�(U��{q�gӴ���2��>G��DJ�UfJe�KBΗg����	ʌGL�S��`7�֕aT��+l��	�����S�v������ C� 6N���w�����ZI�ĘR��O׏2�]������c���Z漜j�&��ݳ�'�;�ZV�����acNA"$FBE��o��Q�i}�n���/�w#�J	�Q�?qj�y~�+�V!ɹ���߱P8��8�/�哕s�C%�a�Uv/!GK�{���wzs��m�؈�<�����S���5���5cӈ��0�+���F���Caإ�����I�}�C深ڬt��	�yW��A!KGV����.����`]�rcJ���S$_��B��ѯ�jI���<���_8	�^� �GpB;�����]�Q��|~���L`aǞ|�|���>QS]C��*���g��>�cV� �+�L%~]�T���^����"�荥�Y�����6{g���=vD��)hi�½�2��>Z	�W�wS�(��IV��8C�8������c����q�������H�	�n
uX�ж����j�������qX��5ݎj�3�q��X�ǲ¬��)���&jbPʆ� nz�Z���pĤd�'�Z�K0`\�2�}�0�\��T
Z<��X| E���y��t�!?bol��n���>�W)d��� P��0M�3}���V��c�P�X���ʍGS�.��6�.G���V���)9xT�:�P������&�ˍ̥$��K¿�
r�����:^��=J�����gW���~����'#�ޭ��.��?��%��W�aFD�6(�<y,7���)"֘��ċ�{�:p���6ګ�rN�ըa�^G���t�b������6|��<�O,�%�t:h�t�$���g
4/�����ʣ�b�~S�����Q��:ٺ&�"D�N�'�ʒ�J*8�����̏��Dj�ý˭�' ,���������?��@���8���ql�&���7�濱_�D �(Z�FM �����&�� ���4�j
`�l,sY]���5�b[r����n����%h���Cq��ZWjw�-���7��p�X/�tcڪ���{�~���>��U?���j ^
������X���yrJ,����=�`��M�o����s=���{+����t�b��"2/��65w�{/]I\�V��wΜQ�����E=bLř�Y�E
�����1��n�ۂ�C**�� �.e�A�AW4g��3;Go���F��R窜/�[��_��Nq��"����4/���O�D��0�P�b�����l{F7�[E	�~�Gb�����~������D�0�*��q�֪fE�~x��d��q_<��u��s+��4�z�~��e"/ꄭ����?.��Dx+<����=����(ЀF�4B�ػC+,�ғ���-�J7XBp� �sbά�'X�zdp��p�}l����Sތ���kYeR�sى��	d
9^�d���s8B��9��-����)S�n�ܤ�KmN��l�F]�巶�$�@i�{ъ�|�'����'�)$1��m�HL���	��h�Y��o���Y�VT`��_�W��c�Ŧ��P0��J?�agNc�hfg�@ή�b���\]R�������֨��m+�V��Ō�1S���3�1�3�����/TI�)+|K;�^�gf�s����>;+c�L k��S���Mưk6��ח9/�IIIb�Z�.VS؞�_��ˋSih'�2S���%��ښ�O��ib1}�[t��P���ZB���Ӿ�>mĦ,��*���v`q��M8���c�a1�c�̩���S�F;����L�@rٺ�f�X�21=�iq�\:@"�׭"ߕ��˾�h��B?j(V1�,����Ƴi-�TF�y�Hӗ
H�F�S�yK�!Y�!e�y����l.��~r�{�h,���$��J�t�b��A:oyY!s%[X�T��q�S|!ܼ��=�+� �1a�\y�}�G����Q�Ig���~�X]V�v�&x���r�����E]�����\���|�k8#2\`�M}o���DWAǤ�h��>j(�+7�������o9���C�p�B���h~��	��hv��ЮE�{�^���ӹz��pd�2�>�+����*�݈z_��}Z��]f��~��l��nZ�nj��%:*�s��{�<`,�˯~�t���Y�9fIzD�ޮS��=�eZ�GN�;>�#%eY@yU~f�z���Q聆�p�iB��cLTT�1�%��$�w!��]aЈ��.{!H��]�_�#���)WK��,�
pɎ�BJ�&U��<!��˕�ˠ�R�ԚEx`���[�b���gq����ذN��������jC�@�����L�c`p�s}�����c?��t�4�0Hp��*�#"*�Ӧlg�������ۋ˭����!����e�b�XJt����\]&Br��	ظf�[��]f����^��u#R��Y�1�X��/A�<�t�V5/�+���bܼ��kэ�,ї^�lS��rV퀄� 5��j��v��i��L����o$�ln�Yo�5c��I}��5��������2�V������@
`	^��$3��@���	n"�Z��������<�Py�t� R: ���0��>�HO�+��Uig'�? ��Q�b�,���mC'�0����]:�����w_(Mv�LC�u�\�,"0��f W�@��҅T�
�j�{��0�{a0(=�\����:�o�yw4��wϋ,��`@f�f'$��VU�.ha���)��\3wٸ����,:q1�#3�gS�_��7�����`��8�����F���j�m��)��LCX����ew~�?�J�k+�m!x�m��� o�+�d��ッ��Ȍ �Ų��!9ސ�����Y7�@\s�ij'H	~����@�~"&ܞ���x��so�1_3�`�\�δ?ɉ��4�qZ�LU�����g��֞�#�w��b�_���"BD��	�R� ��0����84n�^z;sV���B������<��<=S��'�૥썿}A���:�Y�"TylY_3�<q�M^g�2v�[���>�`U��Wƺ����˵������r]yN�!ӂ�~��,���쪴��utq`w��YJ�z[��6�V��Ձ�4N�#�����e��3t#��ec�9=M��C58�1p��Q,�ɀ���[��c|��~Oz2f�YUЯ/���o�Rj�O���|V.b�ba��4q�3��&��f|���i����x^{lyI��n�G��~��JL�p��2儏]䐵�!�ʆ������;�������E�g�`�@�����	�hF��8��6y;?��R��Y�]M�oW@���Wq�7U@���+��.-����C�-`�i�0�}��Y�Ù��xK��>������%t��鐚��C��
N�~��vN��\�~��
��!6�۸˚ =�U;q��)��7���P�T������ɸ;g�e��D�fVƺĸ]�~^N�A���i�ư���u��|��;�-[��|UK�#ٓ�o�6A��5OZ4��}���o�2X��r�vG/�TV��f��9��2q?�~��؟?�-ahb�|lx���y|n����Re�ߵ�p������e&�l�WBז�y�o�$��80�ͩr���l�+�A:+=-�������<��>تp���P������ph�_퓁,��l�]dBY���G|�������+��Z�p����޸"�8=�>��_���2��3�E#֒���
����?#˜Ypz�H���j}q{c�jL�:�`W�2_5K� m������4��N�_����d���vZ?��:<�4�1���:��x~V[ԉ�:�I�����Eϋ�w�z;����M��Ax߽q��!6�=_��
����C�h�+.T{�ٻn���~JC]�˼m�L�����K�8�&9�f��0�W� �S����N{ׇ���y���������n��um���LoW�<dQ���{>�FH�0�=˴�������Zn^����C�ތf�|`8{� MY�������&�l����y/%?x��t>���V^�m��l�a��nz"��8���rn%#]�s��#s�ϵ�n���g�Ԥ��9R�@L��FM��P���9��QĀ�SD�L��E�����4��Wd�9�?�1,{L��
��U�-�GsQ[��xV�1�kE��%���]\^J1�M�*8��QT�$<q�0��w��4:YaS&ه|vܞ|J\#�rB��3�|���)�l�
�R�/G�T�����	=4�scd�*倶��o�xi���vO�8i���Ν��pR1��7>�<��uWAخbL�i�h��ȡ��&��n+�E����S8^
���e6�e����P�|J-0K
sk�"r�2;9*.}�����B��{2���7�wp�.E��h|9�������u�|���7�C_\��:�Ǜ8���ArF�<�m	�n<� �Q�n���\ m�e�\���!�w.$3�|R_�*��(����S2���d��������i�;�@	&���O#C���g#��v=��[�@&�?��`��ܛt#��Rxߏ���?3�7�J�U]��C�?�پ̚�fA�a�3���n �?��O~�~7t���~R�z������~ʸ���(�+��(5����A��u�?�EQJY��0��]���z?���>L��TH��k<�J��/i�҈�')Q{P����p���x-P�5��Ы�Y����d�ꋚd~^7YBW5
\��U}u�ڲw����E-�&wi��G��}��(8'=r����Z@ǀ���t�_�Q7����rf�bny5�X����@+]!�����#mG2�t�{N$�`%�g7�E�S�T�^�:5T����1g�?0���3��d���;E>o9�8Ԡ�z�&RU�݅EE&K�FkO�K����5E�k-�%9���pf���ϻۯ��r�q�.9�0v�a��[4Δ6Jy}U��O`׭f��h@9�,z���հ�<e�&�`]/]N=ܢ�"[�!$�窒?����gXZ�Cvz�'ؽ�l�#L�Oc�>�&�jY"�lo9.�$����c?|�>�iu�7�?�����{�G1��/�PQ����f�<kb{�XyS�?$�KҜwg��$�z�R�TWU��끺��x-Q\n.����8T	�~�e�������2ԫ���,�(�e�i�_tFj�@�ɷC������?������Pz��D@�H| 5E�t�½��[�S��!�lܞT0#�.�?��T���]bs����g�y���GWC�R�eRϮ`pދ����� py{n0�����v�I��X�2F��XjHJ:5U$��}Uq؋D*BJ���E�EH������&a6<ٿ�@KA�8G �^�n;S�tcdG�j(�͚ZW�ڙKmU��S�Ӿ��m�W~��t;�N��	��((��o�����f�:L�QZ��jw]�u3�8�#&�A|�Vl��ι�	���Vj������,W��	)�y"����z��( �uߚ���a�I�n`4Ϯ�s3�����N�A� ��QgK����@p¹����&��uo��Ͽ~Xزol'���=~���o�,n_�%�v��nh�l���R3�kW�F2#��K�MW���Y�����dp�)ofo����;S}�� @^D}k2ǗW�D����Ӂ��}�/qX��_\9ؓͻK������,_�/�\y~�+l�>�����$����$(���淑ѴJbq*-���4�ˇ���wK8N=Vҕ��BN� ��=���D
�)i�� ��R3��2z ޺��jCC���Z����
��o�1K�~�'4�
�j>^��Ux1*��*��_�c�-2�ژ:������iWme�syvB�'�|Q*$�[��m����bB������a�.�e2��p�v%�ʁ$�����pySg��o\��8���T�����>�O�Q�_���Q�}������9h�O��=�X���<��{�_���vK(}�1�bg�W�~�G�)s������{Kw�&��Ҡ<�G=�4�B����(j��
����{2,{�o��t��txUD�p��
�a�;8|+
rg2��[^��|HԞ`N���?�'���#q���Ic;�s�	e帡1Y*F���H6�֡����������Aםʐ=i��Ř�34�2Oހ���IǑ�#��(B8S~�thT�^�Q�y�8Y[��9`0��'T��.)?{JوS+� x^������_)�6.�Ra2l|���Z|״{�N
��]K�x3s���|{9٬������km,U��f~Z�+`=�&�K�8h�WS;5$�p��:8�'�&@h:���u�?-�l5^XX;��]�`���P(.�6?���	��!�����I�ֻ%r��.\=*����0g3��\p-d�����o$�&��\����Tv�>���O�z��MPU��QTS���.���Q���;
UV8ׂ��Uh���f�:Sm�&l{q���Bkpѱ����	A<$(�:�ϑ&M�e���`�O։�J��!&bj׫%�V�t�P����{��x0"1���t�Z2��G�3s�=����k���4�h���Z���~�Б��!#Fz|ۨ���VV��AH�����Վ�,$2W7�z�X�R���J�8�
"�W�D��3�<��o���Yh��G���O�Ϟ,l餸5\GF3U�d�$ܙ�s��:6��<�u�kA��{�f�!��"S����s/vf�GU�K��Sy��+��}�R�H�����݁��ۯ&�����`�<2k�y�r��P�q�zY�����:�V��ܚ�\3���|��HkBk���ʀ�t!��/Y�eZI��si��/��Ù�tq�����e����?�ǝ�������ҁR���sV6���UóH �t����;�eeg��K2l���w��IA��>n"ׂ�ȭ�6D��������e�:�n�?��B���~]�Ҿt�I?��(A��sm�h;�J����]se�o�>�NÃ�&�(t�L��c�}?
XV'	uiCXX�\X?S�hp��e�Hh���Nۆ�F�����T��AA��T���Wް'U���m\�C���gJ��}���΄�����C��������Z~P�:HX����>.�ü��'��}��4s���}C<(�\EQ�	%���O��,�&�Ev��hb�}���%K�v]�>!������|�-�nb���7�M�T		M+��>.oK�4���oe�%l�G:̛�ai�;A�D��۟�"Ix]�#&���ÆC�8%3����I/�!�s��k��WU��Q;}ti�Z8:�ω�V[�
�/{#L�n���6Oк�{�{�=0��2�fb���Y��a��?Fw���oL�#�/�X��ֹ9�l>��p���ۈ��%X�� ˯�R<�l������XfK��������/�p([�W2I<8F�2�>
��s[4VK�$�Qӥ@�t��fS;0WJ�W���$�R+��.�
�\0""����H�k�6���ө��Y���~`�7::J(hձN2L��� 伹o���M�#v�v��ږ��(��E������̤��߹��cힲ�Rox�
����w�@1ﾟ���k�0zA����:�(k^����ٙy�\r� Fq=�u�co�c(zv_��Ƴ���ǳFW��7x 
&˸��{zZDn��	H�����e�'�r�tv?\?T�y����&���Q7�a�+_}[����������g��g����:�I$��΋Xǳc�W����ā���G��w���/�;�xOd�?�q�6+|1�e�cЦ�!Gp0�����#52cC��W��W�@�� �����pQ����m:�˒�E$�Կ��D��� �p��۶R�M	��0����6+J�NAQ��I��c	�'���m��i=Gs,WJ�΄jAv'�4搕

+a��$N������y#�5�,Uձ�~R$��}�ڷ�@U�ݹUgg�Mn}8[���D(�#B�&�-qo+o�C5�A`�,C�*�t~-�12"0r�/h���~hS�R}�z'�tƩϗ~��[��wOկW/ޑ�v<��$)�.�P��u��'�4��8fGP�����0=��b��!�X��Zrѵ	��ZX#b5Č���ݤYԤ� \�u�y�t��r�`s]�{[]T�u��Ÿ�Q�m��7���6���H��|'�����m�v��E�n�_�LV.��F���_�)j�k_��gQ���{O��:+��׼�L���Ce1��3j��þB<I�ۜR�4\Q@�Z�gӗ�<i��}|��Щ��9��B�Y��� ��u���xZ�영�Ö������/��ި�|��Yn��sea&�O}#�V�#4�L��w���jc$bҹ!�Oೝ0���5(�Z�]�t.���E��E�^s��K �s�i'ô�&A�v}Lnf�mF�nD.�M�E��EX4�Z�w�G{�ic��=HfƂa���ns���.�l�����d>ʀȏ�]��L�YyQ���u%�����\�@ӧ��Ern���|���d�Y�!���'2��k��\���Kw
2����rA�ֵ�s�r���aS�s�� �V�1��$�b��Ͽ2�6���e�jG��p�#U�ƨ��WK�Tp7���ܜז�k���a7�t7lO����,7��Xc�j�!�D���͌�zс��Й:�oڈ�V�%�7'l��Y�xm��SvD9��Mn��ȱ1��ꝬZ�>�M7{m�ʏ���K17��#��'��XU�,����=� ��E�mI�DM9���^�Ӷ���G�����.Cۣ��������`{��+��S����s^�&��\92 ��(x5�`c}�����u����?�b�,����P�F�F�u+8����y����
4.�X8P���S��'K�s~���k+S��Q�kN�o��St���>0h�����9����L�|�sӍ�"aV��yJp�+�\^�P�a9}����7�d���4%xD 0+a��*~Gq`���I'���Ok#���90_���m/E��ׅt�$�`4���#q#p(�uѻ*7K��6{8��7�#��aL3��{m�V���i��S��:B� &NH���~��^�7��44���A?��[�T�¾��Q�#��ViSF�)�Sa V�b(B*"�I�˛~j�'�TDiA��	��]�a{�-�q�?�QH��.�j'[���D�������0K��R_��I5�$â��>)�t�i
X't؊Яj�N�r+�j3���{�wuD=?��1��l�itw���eƼ���i�.�~�Zv��;#��`�yƽ=�ōȕ
Ld��$C�@��8��>\�����v?<*ٻ��XZL�F'��W�*����|@�|@�2�O*�N��)�)�X�n��%g�kuC���>�r���NAr�3'Y�u�\��t�P���r�M[$�6O�#�?5�񟶦��l���T��TTzL*��~�5��./1_ sw�8�(����qZ����!����5'̣���7:y����<%�sz�}�)��C0LCs����Ƈ$7�ݍ�"��h��S��W��ʤ�����c��>~DcrH�n�]�6��s����e���G��M��G�"|P���f��v���+{�¡"�
C�cm.g�>�9N��u4_g�v���l�Fs|G�6�X��54H���@IP�a�]�[�@�Զ��|;~`���y�@�To	챰C�噲�&A��KY������rN�AX[Y��U���:�K.��2���mHR8ێI1T*I~)r.���� ٤�q�3�z��6������a��Ő�3�Jb���'��0=�߁��v���1���wM+<�C#dw+����l�_�G__��_���ӲI	��V;��{�z`�?�1i������ʋ<��C?��|`��E�Э�û
&F�5���.L/;��B��&���X�+��ْ����ٹ{�uט0�Hw�#�e�=9gwi>�6�tR>�����9AS���"����|bb�H����$K�θe\2�( �M�/���)�zΤ�����\dHo4ѼXȿڑ�Ĭ�/���W�PQ.�������h�����݄>6���-��s�/���a�ˢ��� A�{{��5u������tä�� b�ř�~r�N��|�*c�z�$jE�`f�5�	2�#��ڴ8�~�%��PW��]F#q��H�{Ѝ(Ny.]�M�VV��*$z��v!���8��h���n�mG]��]gd7L*�����U�%J]�T�{^����I�Je���-.	�	�V��E���_��-�M����R���嫶���De�3h-��3�bt�Bykn�a<��A��+t�Tۃd��~m��W}-F%�$A�|I߫r���^*n�Uז��T��Yz���CG�sߙ���j
?⡱<�|x	�h����*�#}E�|-&(΢dk�t�۴�^ZX�O;�@-v���ʗ������C���'I�OfZXC�?m�y�w.D%��c�A�t!4O�*�%WW������!��;f/}��Is�D�>А$�&�1�蹚�:[��&����<���M�q�_��b�$qLIE�p����b����}���o$s��x���_k����D�^��TUf��J�R�\�`E��s>{� y��mf��4��J�~g��3O�yߑ<�DI�D=��TGa��<笴l��u�Z����HH��E�Z��2Xo��ȋ2�9�˱����T��7�n7bW�m�S?�K�:dD<��[�[�'�:<���Wl�]�^8��ײ=�q����	�p=�YА���9Q�,�nw��N��w@��U{_E�l�]C�)?�}{��SƘ�zB�Jyq;�m%���s�{q����u�css���]v���s�q�<>͂m:r�/��c��k�
������v;J���.+e���+�d��9;rl��Q�.��֜��+���e,.t%Xvm��f��ZŘ⌨������f�D�vcꈲR�SM��H���yKf��ܦ�'��)ͧ��C۵e#	�EX���b�Dp��r���mOr�&��<I����9s ��qsaVuN��݊yOXzu=�x2�VݻS^r�1�q6���Ĺ�e��cn}�8KN�e"ԫ4�J�af��i���hΜssQ��]���Q�"��S�W���Qޙ^��7LWU��ts��V�Z����F���;���M���E�[�ŵ[��!Xp���C�p���.���� �5H��Π���-̠�s������3��wU���U�k�r΋�ȺO?��J�#�d%{-5�f����N���߮���1�aMلf�:���;/��o��X���	�N�X�����}�ORM��Q�4yE��yq���h^$�����ŹY�����|[�*�MWA3ovڪ�r���z`rO<��[aD1dfY��H�<(@!�hd)��Rv�:#�\q0t7iFC����IZ����x��;�$�4(�mn$�ߢ��&��墂E����N���K8�3��Lw{rA�'���L���rS
5�_r���&_����l�
��#�x���%���q�6u+����,���"��@��o�:�7}�_T]ot�k׽��a�k�tlM�����)�y���[c(�͙1�u#���oǆ�IH5�,k���;��ֱ���Yp��v4nog��'N_Ul�έy�~ʞ_pMBt{���IK�z����3K�O`�Ű��S1��[�x[0��|�Beb����i���r�if�kޘz�R���W�lb�<��ป�Κ��44�0ojՈ������'�',Ҿ;j�M�D�C;LvF���}�f,���>D�y��j�����������m �˶Q��3..�,L��_G]owq��7AZ�����I�o|�_c��L����8��â�f\��q����X��f����_�����nU���^�$ɫ>�������<��q�A��''��o��f�I�?���jpkM�(�$��b�H�m��^=��^{���Qz
�����5��F�.K�#(����,��x	��9G! �0�����;a ^���,�3~&�*G�˟>:,���9�#3�Yg�o��k��¹�>��Ɵ�����v����q��'T�N�v�ߔ:@�'П��@��~n�.����f�LЋm5{�]���AhƢ�O	������8�_1��r�tu̘�}�r��I�ځ�Ae	����K��avc_�;_����̕��۲J�u�z�ϵ��u #����OWP�q�-Oh?odI���H�h��B�	$:�E�Ͱ�� ��6��ޟ`�W'��Q� �5����2���8�?�{�{r�.�?'�i��yy��OF��;���	�Qب�=�X��7p������s1رO�3Y�ϼ���1F��
���a��L�к���[��=FG1y��U��\���e�=Ǐ8�­�������|����ʺ�T`�N��[sj����խ�A������M�ry���Y�"zݡ`�ڰC>qR��a���U�')�D��X��Ԥ�����0�j�C��V�>�k��ӈ�o���k>���:r�]�3/2ƮM��� ���C�7r�颊�ʭM��TSk3�ӎ_�?"�=ϋaMW.�"��L�SMc! nn8�"���B�����A-�׳�`ȵ����~;rn�ݸ�
�ε��Y�y>���r���g��4Ta̗L�.Hx���-�x+;NŇr\�S̼���ۭ���:U�������X�=�)>$s�kq^Os���&<H��1}Q�n(�l'���\����fSk����k���~@>=�9����z�#T��ۤ�� �^%a�os:��U�;e�F���y�>������2���e��R/��?�a��UE�9�S�R��V^�����X���l+�ڶV5����X	ge�N/�����+BS��Yl|�a�� 7�*� Z#�1\j!<�x6^���)��)CU����� �D��,��7�l!�^�����S{\��RڔV��~��Ƥ�FDoI�m����0��Z3}�Lz5'b�Ny��0V�3=�o8�*(����b_��z#��!�ja%ȅ)��G�X� Ҫz,1����\�?l}E�hl���U����W7R�2h K�SDv/nM�F���s/�1)ӽc~)��$�@Fm_����%����k)v�o��Ը��lvQ�_(zj���*�R�#����%g_�|�s�SM��^+����� �7���kO���u)��=�/3A�8�.������	3?�l����V�S/'�f����-�bI��lᵱ�<�Uܶ
��U�(�0=QC��c���,�D,U9F�h?��p�`i#p�Z�ZK��Rm�X�����%1zn���� ͚����(��w>�	�w��2��W]x��ФH��}���O��&���M,$�����&�+I���+�+�������`���K�țBG}��U��%�CO����̀�J{��� �F�ٛ��ؑY6�������'?[[����N�~�̉�{� jv�OLJ
~X�9=�B����;r��ʧ"����jN�Z�P���gY5T��O�갣t��H��آ������S���-�M�V~\��ޘO���X#{�l��q����P���5��j���F7+�o[8c��Pq{7�8Y�v�w����#�-����:F������ʐ���3��O�b=(n`<�Mq�J�ܓ��w��z��:�����!aS#KQ�9�5��!^ 9��ǈk;���CȄ���
XN��U�
�`�I�yBG�bnoO�~H�N�7B�X��&���AR3�"z�����N�1�.��4��9W�}W ��qz��3N��v1��u�5������I���\c�g�zu8��n��{
O�Ճ�?���������l���d����i� �',ʊ��S�ɼ���2Q�.l���=��4?n�D9�P�R��`4J�uǶ��\k����d�U7��X�0[����W��,�kh�7׷����27I��@ 裃?3`��Yè�g][]��<����\,F��F������H��IAW	�H��3�a���
��S�����2Y,9�����[��<=��F������J6Ǯ�/��5�������oy��X�|�j�ćbx���"Y@�a�1[�A�N�-t��/Z)��jp�;��L�^��c���0�e���u�����>������mI�d..�؊��E! �ƫ�B��AY� eiH������2F��c� }b��in�'m&�~AM���+.r����Ɩ����}��Xٌ�UP�"��ױ,���{���d�Nh�}`'���/�����6L��,E����k_RJ��U�5=jMY.l�X3h�L���nOְ���Z��;d�w������u��m�;���9�[o��n�Wƥ��5f�����*���D��e-h#�|���0��T6e�¿H�)\��,��l���7�Z��5��I�.��n�4!X��➊5�l�6\�z�R%���/�K�""�s�β�!�?���B�{c���o��X9)ѐe���;仛��{��U���\�n�f���ŕ��Ԇ#/�P��Q�Η��񞀊լ,O QR7O�c�ZZ�����������k�4F��7�w�\��V$x���z��Xއ�D
vb��씝g*D�]#���1�e�7/�=u)� ٨�۪ZQ���`Z����JE�=�E?�P���L\C�[C��*}
Lݏl����2l3�Lv��]Tǘ�����ZW+�����ڌ[����8L;y�qE��B���އ��-χ��kDm��PVY�;�'��`P^����D6�	j��節�D��RˍZf@���o��O���aO��:�7�ޡ��Mhk�D����hd�.:1t�/�F##����x������О\_�J��(
Y@{��$��q�*Y7HF�s~�M�)�X��J6��[���5�a���yJ�1��" �`���ň+��n.����zJ�ΰ�F^��c�F=�x�J��>��*d�>O�Ӳ�����B�Ȼc����{y�#sX`��h���SC{b��}��Z��V%�2�W�^Zo�ү���#�ȁ�U���$�߮wk�mw-4��3Xw�~���|w��VF~~Z��%G ����H��A	XC�l��i�U����������v����2���Z��A^��fL��9S(���#�	/yXz���B��Y��*�H�)��p�̫�3,���_H��x<�_���/����|��LD���L)\�Lfx�^�j7�B�n�<"(d�^őq6YݟN���>��s~:�g��fb��h�9D���L�5�H]]V��2���2
�ȥ��8FtH�!�2�6����f�o~@��ޭ� U-M��3x����o!�EN����ܵ��\5΋-0Ή9�H˅7Ї�.XF������e6`��CF�ŷ�!qM5�F`��#0���	��n"be`E8={�g��d$����	�\v���#o�Zqڥ��'���[�97F4�V�����0r���Ot�`������Wz�{�N9�$�$�q�py9¡�	��H��#��׮ĖH�A���@�ƫץC�m�+݁4���LϦ=�LV�Gs�(�XO�ބ�W6;m�&���{ �|j#������'�` 8��: _��5F���ъh�M��'��/�2���#/�_���Y#dn���ı�!�HU�)|��:�V��n�����7�n<����U�-2wAK�VV��W�zu�;-����z=��q�A�}Nrc����p�zp櫪�zx����t},,Q�'�bih�\b��_Μ{�6?��<?e?]�{S��;]3Od|.�;�H5���mj�S���l�WY� O����m�+�"�M����ⵅ���^ЃY.<��$�@4!�D��f)_�p ��o����XLjt��Hִ�ڴG�六��Mf�t�����.�k2YQ\b�	>�Hތ�,L�/�D�v�G.��>S���+����%��2�c���r�����R��B���,w��|���'��oj��Q��F���&i��yt{c��DVmeO��n�Q��dV�L�yv_�NĞ*�1%g�.� ����1WP�/�֒�j����Z�o��jg����|��x��������ㄭ�U�(�c8�f���؋���scë)��.�
>��4���j��3yt��4�F��m��0�6,U�$�>��E�_/�B�w2��6�!H��9��䟞��k��F�ȉ?�}I�zf7�$g���<,���t��DN���4��Ii9.P2L1PRf�:^��;-���l�]�]m{�]~@��1��.�ue4�7�H<� p���ڔ��g�񦺍�WJ뮓5?�|Wy�F@s�\����E˃w�lB��A�iR��]���h�xXU��W����?uj�d�Se*�j18a��������7U�9�ɵ������M�kYd I��r��h-{�S=�%��=�@��������۶��<�P���b�T���W��(����x��T5^���.@�%D.Ÿ�\j�5>_T�w��4���}��������<ڗ�\+C7vl����cAi>��}F�D���T��>J刼F�1� �<�jы-iG���X�ꩣ��y����9\��c\�+��; �sMS�iS��. �S�&G�h)��[|�����z�Ǹ�u��1����5ԧ)����o#��5��K!ޮ4T��%f���k�5.2����nL3��X3� ��A�9W�)��Z�k�K2-6�����l���80b��|k��+G4��GJr�K���xq����f��I�I��5tܸ��P&`M������bs��:^��{��KN���t����Gq����I�TIP����#�n<��16@wd=<G�7��Ÿ�5HCs���ݭ&�C���X�����掼���`e��1D��*�������O�l�l���.�`��9��CD��k���6:שC7� ρ�D�5��x��9���h�L��{;B��*M�"���X^�G��+�ȷ=o���S�+�6��Q�dq��p9�"*v���#O3�:D���kB���Z[�.�9�?)�p,3i���:D�:���Xw����^sX<�lK�iMJ/�=�$4�4��D�����$��{� k6�t٧,�����ttls�0b~;�&��EY�d	�S.�堲q�3���N�C�#�/��o�w�	ߝ���ț�X˺�Όx�qu[�"kf�u`�ֻ���cb��_F����I�o�խ����

ut�^UE.m��|�׻U��_<WT�Rw�ݸޗ��V��^绮N6�c�q,�����YV~��H7�\�����k���'��bK��º��~��@��O7`h[='�cUf|<�{�:l�x�E�fmD	����������E���K!'�5�^ڻ�PDSAÏ#�Bi�i������c�]��`6xѵI���2��'�n~Y��u���VU悬�����D�#؅�Y�,���']��rW�o�<l/$�S��3�|�)��i�O%�z*�;5X���,���}�]�K�~��z����b�����	�Jwx9@��II�E'��ˤ��,���+�S��ϟ�Ak��ם�����Þ̟����窠)��r6�g����	q0�b�� o{X5��tqڏ�w}ZE��i0;$�|����Uv�
�!��冎��?����m�s���!��9����#������Ug��m_�䝜�Xד)�;
�pY��a-��|���u94�^m_{�{�қ�:u�4_��Azd�����w�Q�>��^�A9�[S��K#h�B�{��I�r?}��5��H���<z��.f#ƚ��[��{��9���O�b�7k\Z��N�cs2iR�n�x���4��$�ʼ��+�s�\\�F�{�b�,�Y��0�ݺ����6��*�X2�Dv�ji�7�x�yX�!�wU�9!@?"R"���&xWoo��^��^��K\0�=�ƌf*��ȵݽ�1i�i��E8�j��5+�-��>��"�@���!�V���1f�I�Ɩ�6���y�/sQn�*W���=2��]5���>8#3��!I'>�=)/a5�5w�;Tr��Ԫ��?j
����X
M/!�sqA2�X�g�|)��#��NU�ewq����{O�L���Fg.�&P���W�F?�����esNB�y�����'5
Dj��!<�&�#����|Ѱ���)E�ى�,F�tt�c���8 o;�a��HR�7v�v�xB92_��u�N����� ��O{�k,��z=���ƾ�)�����d�E����Q�2��.�l^�q��5�����b��U��>#4�Ԓ�8���t�AӀ��,�Ϙ6V�:d�,�R_#�@�5�F��|�w�����]S��3��9���Ĺ~�_�a���ԏ5��su{�p�}Vr:��q�?i%�u�r��'6D7C�����I�����\e���2��}BEO�q`������;(�Z<��C!/�Y��w|�������d�4�U���e,숂^KgM4	�g.Úԁ��8U-q�����,r`(M�g�:a�f�A%����������:W�M�̭;8�� �H�|G>��8��%\)�4w��ꡎN2��Q̨nS�Op0����dT�EjB+��%Q��s�����{��h{�Α�>�E�nS{Tze�-���*l:�A�F02j&��WCǊ#��)�ߠ_Z>y2�F�Oa�b����\��T^+@��G�SOv�z�}i�܉?�9)�=L�5���׀"��v"�d�W��s�Jg6P���bR��y��}hy*�v���{���D���l�so����^�,�����dɲ\]��A*�$i"ʗ%(i�9�q�3��>H���FK6m��?�g��"_��i;�=E�����$��_V�R	���;����Pɖ����V��n�~
R@��Pc d�[�%���(��?	U�ݕ LH`ꟁ+��sgv�j�Ȃ:>�Y1���mom����q8IP���;sV,X��k,�8�%( �=�ZM�i�����stb���4�B5Z0.YV�:��+�ă�Ĝ��fܑ�����rb>���Gܡva �D����j��v� .�q"+ד�|��(	Y���fp̾qi���lQ]��y��IS��ǯ��ӗ�n�:����w��bԚ����	�����EK�ϙ����wl�1yf߹x�q���mK�v�M���'�t��x��ҟ�e{��j��!�|��IJ�g2�O�ݛ���	�u��"�˲��MAA�E��|��?�_h� �L���vԻ����e"���*���!m����P��]�Q�⥈Î��ґ��'"9���]�RS^%�������5�~�y�l-=�,���'D���+_��D2`�~����Z!m��k�H�$`�U�
��}	#��T��P���ǀO	�o{��WF+�\&EFC�K���E��᝕k�~�M�Un~7�O#�VaO�G�w>�>؅"�}�{L�v��s
C�֧���a�>(�t�Mվ�@C�(8>P��S�]�l��A�x+޳��d��^]�qp��Y�dix�$y���Y��cl�ΰa�Tʟ�fIU����P64�D^��)�6ɩ��	�2�z(A�%��2nM�XYo��+ʭ�5`�Ǳ�1D]J��}�>V>��"�Q�πn���U�B�Q�0�㰹V%߻�xbt���˓6��Y+�9���5�h����6�$��9S�'
�l����qj��vf���zt۳:Rze��dc��C��M[����������i�;O���>U��/~����s�j���`���#��S����w����������M�zI��gz�ɂ��IX��hk����A���l�)�(�}X�}A�T~ǳ�W�/��6��:�S��!3eIC������Q����q���8��x�/|�/��[M�D^F�10���P�R�2�f��s[Q�_� I��"T�t��/�$\ᖌ��y\�C�\�]�T��U��������,�Ə3��,E����z s���e���k�&��k����=��<f}��>�tM����J��fm;���*[���BH�&����c��R!��"�lX�*�TSd�{Q�Hn�>����Zw��
�u�w�v3���m��Ÿ!��l���^K��K�,3^�	�Cq�!16��w��N����Oo�p�'H���s�HbYX���֡��o���D��4���R�Xg<,�yYK�J�f$t��#�&g�u����WN�r$�]X�NM߫�.�S�E&Z��E��0�Gǖ�W9�@���Ʋ�'Yv� ]����p��W��U3cgi�����eHz��"[�a;���on���L�G]ګ�~�eg��%w�(}��ڇvL=>xPƽ�!q�\�Б�ު>gH�$��V9�c����х�F����t9OAnr4���	R1̌q�M�^��T\�̺ʩa-�z��[�N����0��΄���Ib�=o�g���=��K�j�����)���Y�z���v���@�������T3/��⟂�F�~3���t�W�G�9v:bC�����k'�r�X�tF�l�����CWo�W�8�KI��zKL��!�T��qL���,�"گ<}����6�6	�6N�[��Y�9D��k����V=7�=�pmC��������l.<�AXȍ�1SU&�`�FR�V6������n#[�M�C�i�:F�j������V��=�?�8�vkRhK$�8I�#��,u�P�%��ҁ���u=���Q �� �x
����wg�qs�����H/��n��^�rM�����;n�:\$�jG�(:RW�xG��si!7��B��w�Zuq�-F7Ne���ЍMv�}� ʐϐ�6�o$��w�1,v�M<�+�$�m�H��>G7a����x��!Ԕ����E�ɧ��9I	K����:\8'Z�q�}5p͑��r+�}�t�����H[�@3=ٟ��yTP�M�˝���M��)<��
[}ڥ��Ź��=�;�!�r����*d������J�1�F�)�a��	�k��e�CbY��)� �7�h�z��-C��p�4�-6����J�}�N W.'�����큱��|mEw;.,)�{ �Y���#������ܔ��� ���nl:�P�1K?3�Gg��>as��������h�h���a�H{��X@X	cC�9�Sv��)f��G�!�N��?�o���#q�uϭT����&eb]�t�`�C"vfa�ʬ��r�(ہC(���S"���]؄���J�_�p�Un[,C)�(��#{����^=�zC��c1���J��T��ᕏ���;v�����ULGG����c�K�t���������̷o��F��b�N����Dk�Y'��m�'Ry����ƀf���}z<�8�y3Ή6�y��Z��6��G,�r��Y+g�
��\�٣C�VR-뺌�#t�0���}����U�j��\�yUy���O=���7f��:�*W�(�-K�1���Ǹ�1:t�;F9&T7M���@@�Ax$�T@.�3�mCu�Es2�
���`�1�c�;��1cS�%V��>�#�]�kN�q����T��ܰ��I:nva՚^�5)�>$|n�Z�����za~
y��٦uī�UO�� ����^����zOq�Ȋ��K���M�8ipF��f���{�����*����bB���3#NbSq�5+c�I�l>|�|�&(��$^6�y1^�Q�)���Dńԩ��� �'᫇��Lސ�DӪ��]��J����!��3R�1�&��R�z�q��ב�R�(���|�e�tn)h.�����7�f@�>��)E�3@Ų��Q/ '�2�o��I��1zi��������#U���2�����id]!]����fO��VZ��A��sS�D����ʧG9l��\|�=2�ƍ��)A�c����1=cV��߹\
�����x��	�A{�<�4�|AJ�o����#7��{u�!w�!G\B�c�;���~������-�w��_5&m�U�{x`+�[��Pss�G�l'�;�,���F@�&����u[ڑ�b�'�~�C$����.FP���e�a�W&���ȋ�N!��m�g ֑�<���sK0+2քJ��r�|��z��/�6iݝ`h�҆�����S�I�g�B�u�h%@��o�E���Smn��&EW�|�R/��5����oq"V��(�O)H�\�{�)#�׆ƈZ��lݞ<6Q�S�ͻ��}ĄW_U�|-���b�?ͯ�&����.���TrJg?ՐVA8���B��`�sl�6�zѸo ]3�p�LV פ�)W�]�@�V�g�â����EA��M�a$����"�'�&��r{�$��w�"�|3Ak���K_��"ge��*��Ŗ�������Xۏ䶤��&ɛy�f5�͐|KAi�G!j��q*�.;���������ieUe{>�;���	��[��ٽ��WqJḭ�C;P��	���V�E3�w�Q=�R�bq�Ջpg��J5be=���I�O[�ꔔ���w�2���^�0p�rw�7#._O'ј��"����
SUzx���*��!MUm8�ފF}l37��i�Vj�����^_���d~;�3�%4{;�g-e+i��RO$YPA3ȋ����XkJ��g�^�aQ�J$��tt���Fk��&8P���27��5�xU}���:��þئ��Э(n���T���1u�nc�٩�p�9���D�>���\0f��+{��+	bGA���+Y�6uюo��$�h����ۈbD|=d�~���g��8^�?X0@����[c�qI�i��G��t�u��(�s;X���~˂͖G�~�������c��ͤ�6�ށ��v��1`��0\�|Ň��[��
X1�x-��z�ߓ�n�r����j�{��0gRJNwE�~��-lhj9��j�Zu��(��	��*v��bi� ӥ����Q��K�|P�4[/�9���|��i�v�U�Cڇ�$��:���<p�Q��.[C�4�CskӃ !�h�$R�3C���SWթ^�j��O�)3!�(g$]f����V?q<�ѣ��D[�pB��^p#@yp$�꾁�%F!�m�,5��e��1Z��Qf�)(O􀤫��*��f���ӗ>���8��Td��7�Vˤ@+yΤ���m��@���9���=<n&z�ug2BN�KO�?tW?	i�܂���̫�WJ�9|CĊ� � �?fk��tv5=���QSB�m�_9A����,,�9��(
�\���־�~�T��&�~�g���׸x��|�8�XzU��n[�N�ҍ�S�Ag�JG� ����!��I��B���f�c�$+�#SrnNR�Ƌ-Ј�b���ͬԅ6�h�u�*�>�fsc���䗯�;(��'&���[��R�?��ȷ�\>v��~�l�j����t'x�*r!���uUMR�����W�������L8�]c�F�9izQ|h:�k�{�rW���o�DQOE�2nHϰe�^z���Cr���&�^� �P�SE�`������D1�mgDn�`�:<S��p��f��'�݅&Q����<G��Y�h&�Z����;���%��ض�9�?�j�J0�`/a��fu���U�s>� �L}]��]�oj#���|�a����g�dK1�� |X:���H��֡����ة��Se�o��<�	��Z�N')� }yM�1��N��Ʊ귞;���È�$$�v4��1JWI�?_a���-�"��k�	��uL��{o��`�弶[X����a�&�7�%e�����@N�*	���F\�{:���̙�me�?���(p�lut!��.�)����&3���d��e㧃Q��lN"^S���%�2y8��(W�G��N�G)T���M��2��s�p��_Q��Fc��{�F�d��Du(��VC_N]l��;�����/��ޅ�����go����ע��ݙv�G��P��MZ�^{@�K��Rt����/ ���%(~��w��3��9J���@��<,�NdI!|��K�U��I��m���˜���nh�6���VW�O�o��GT���0�4~?a��'��٪[mk��n�$��c[2�D����������W��,˵��7�ǉO�ݻ-�ߨ�2���x&��/���_G���v�}Erc�����"�W���R@׮O�?oo�	�;��I]�ePSB�ڣxil�|��~�q��:�'~�Ƨ�S���(�n٥�@�"U�k�bB�ԝ�kh���UHڝߚ❍U�� ���c��E=4�C���8��qxs�����h��1���q��.�`���,�bтSG�h]�eLg��ae�潲��+�7���?"1г��CIX����U�Օ[]���=Y�4�Q�f�>S<�|}��c��g���zn��XG7��*�۸�X{ÊnX4�������Z�4��4b=L�Ŋc�O{��k��ԅ��P�,Q>J+����f
 ���T�F�l��$E]TZZ��c��|��]}�{;s��I8yd���5�7�2���2�g2��Ѣzc�̠&'
��d��u�!2�i�״j\t�-�eŶ�oOYAx�48ä�	��&�D�C���ⴱT���_PZ�)�U8aO�#�"Z���U�����Q9�O���_��+ݣ�׋������c�O��V�d��|79����4'�?�W��Kw�8����?H�Fc}�Wtw��b(�pn�O�\W������cܾ�{�y���M`Z�����ѓ�S^��ܦ'	�m[D��7�F��:2K�"�c�;"CYq�/R-��j	R�ݴ�FŎ�T��Q��K�6�e�;�Y��_����H���
�
��	�29�@�W�4�j��s��x��`t��Q�wB��,�����I�_��������~��|�i�#��+����<v�H�Jܧ=��ӕ��}�)q���^ ��j�5�lL_�Z��P����2%%�Ǔ4�.��p`(�D�5w�y|���㱋�q����^a��zsɅ���J;Z[�t	 &��0��V#d�G���b�qjy=P�qh�)���D���	gOp��Mpݿ�UaKM�����KĭρS����e,�����P��'T��-�W+9��f��PS���1R�s+���F�K�癒�#w�_�v��z�/�:��NV���F���|ߔsGI���qm�
�V�i����?�����b���6�0asno~��ʕ4��	�-��K���y�ãk�5��������_�Z��_��5�z�o?��]\�¬��~e���2�5m)Am��x�-�^��߇��%-k������,]��k:���o+z��R59m&f����`-�.�.|�a/�!g�4�k�J�P
e#w�j�緀Ճ
��(kF�A8�9h[/�mq�{gj}�����$�sO^xH���4��͈�RiB������@�wH�'U�VN���N�&����tl�]e��\���w���(��ۖ%��M�]��q'�G�W f� 2�N̹()2��/Y�x�W1�\��f����L|��v��g�0t}�2?x_�	������*���hp��їw9�˥�i���]8U/������7Y���#FؗAl��}�a=C�*���X£�/�K<�e�2U�n�Ƿg���L��O܉��Sl�g��X�ڳyZ���џP��k0@>��p��/�D�i��y���B��5��	���0+����ˇD�e��q�Wf�� �����T>U�����#�۪�'����	Vm����mB:'�P���ǘ�V�ԽY���\E?z�T��u�����^�� >w�<>֡���ެđ���U�7���T_ʖ�<�;%I�0l�P�rǁ�l��DO�Z�>6���{�{7�E|ϸ�jD��Kgب�>T2'�� n��PyL�=����~iD��������em��gR���e�Y@N��YƆ.\�:�˝��������/��N���`���j��A�A�p����������t�c3OժY)�r���躞�g��L@�uLG�>��|w��<(�OXMv?Z�{W+����W*>n���D��S{�*x����e����E3���Yڡpq��o������˶�\���B={���r=��/��$V���H�7
Yg����݊?����]V);�����!W����'�^���1��k�YO�7--t��d��P�V<�"��M�
�R��ɦ�6�-iA�~,!V\BϷ8��!��:��Zf�}���v��l�$:�H_.l���5��{���g`p�0}��~}��)�v�'l��gr��q
�֗\�Ą���D{�4��q����G��e_`�!1� �;,n����[��������4�i�-�U�[�u��)��FT���ϓE颫hĐ��6���}��Aݑ�z�4Uj������ m��^d��jF�&�8�^�m�=4?7�OrF��^ͼŴ#\i1Ͽ��\XX�"m.9�238B�z��6�zs͏rpA�iW��o֋���v諓��WQ�]?%叼�njh��u���#��.g/��^቎GZ�	����A�pp"���q�/�I��� ����q�S=Vg��U�.SW�����yP���;�÷K�6���8��1M@���"z��g��.�W�;'w{�/�v@�5����w�T�c� *�l�>�f;	�,��7F uV����j1W�.BW�ua�
3-穪N�Zf�Ѭ7u�ܰ����ZF��~�����޲����-׋T����&�~����T`
����#>ی1W�����I5�)N���j(`=�
^�&����(�<�3����l�%V����+]�5;'�����v{��_��v.v��Kv��o��	��On���YU�z ^��87�b����>u%��A��$���L�cPz��9��ҽ_���݉��pk�P��g�J$��ؼ@��X�/q��J��ȝ�bZ��_����l�|�f���19�+촴<FH�Pf�'sX�^'\p�����O	��c�I�,���I��ؔ�U��iz�������z��6[ֈ�_mF;2q�pT�,E)��G/��X��뿶�-Wha���VXA�2'y��.U����۠y���7�I8p�Mlq���$��}IjU�9�1b{��F��
��*�(���B�|^�� iŇߪ��})
ӣ?�6
6Ҝ����V_Ig?iP[���>>���tk���*���d�
s���������M�>����+�/<��/0=���v�n&ә���8�ʠ%;�A��"�|b�t�\�R$�bԿY|߆���=��r��_�D_��F�W"��ΐ��_�~�Ԯ+RTL��ob�l#i�����܂;J�}�ŝG|���8�>b�~sZ<�rjԶ5��}�IzY/O�x��$���y;�v��ZH3L��W���5^P8z�ۯ��f���i�f��R^p�_&��Z��[�
""�5���y͓YR�����l����K
_r���R�0��\�Vyw�b��׶W���.���dg���68������4���J�!����jPE��������{xx���z���ڥk8�f�w��tl۶m����ضm�;Λ���9��c��c����j�Y�\c����q�<��dr%gR��d��N�N��/o���h+��0��T���$�5��@sT����z`e%̹��M�����}�m�V�i����d�%I܎d;���j�>^]"p��5S<a�'���e��v�����/};�`�����m�z��#���ю�K'��1��m�Ư{^���+
��ۻF�n�۝�|����a�"��+p�u�)�=$/� gr��=�C��u�8dP�9R/J��O�-j�F���^�}���!8�H�#�h�����M������;����Z&_�Pu".GW�g���%"m�-��8���y,���}c����:Y�|�Ԡ��RjB���waΎ&�T�L����sK'�Uw6Ŏ���h{O�BD(�	�ڸ"��L����A���ت��љ���`Z*K�Jd@�xb4	��jt���1��}�+�4�k���6��3ޅ�t�I���>T���kJs�Az�$Pi�wǆl�����ࡽ�H�+�pǁ���.ч�.rMM
���T�?�\�>����T���g�h��뾱�V��n��x^����O�¹Lh����gn�<vX��^	��T���(���_,��������"��M���񛽽뻿�.��"/��8Ŵx��yE��-�-2ʄ%��R�ʪ<���9۫�ݭ��C�*	�$G��O|����'�
��N�9�"��P�yi���UQ<A��!�2/�����3���I"I��4���[������Y�D�j���P�i	\�Vi���K|
�z���O�����c���_�b��P6@��+�{e��$�525���^��fwݩ�=_��q2��;��
���a�K3��,FJ�iJ���ѭ=_�f�` �p��Tӥ>B#�~w�j٭���_�d���^�q�9���yjg���>��wh�V�Sd����Hߍ4�Nݓ�3��9��Cx���i��w��M&�N�
��Ć�^|\���rҚf� ���8��E�4K1��.���?ZEXyT먍�킀|*��1
���;mR2�y���t�$����3��,�{�����V�f6�H��Câ�[{u�=F:��W����}��&�޸X!Q�.��>J'̇���ui��E�M��Nf2Aٳ/�>y�90���o�Ywe�S���8{�[���5wZ���?LҠ�SL����E�L��k�G�q��;,�H��ie���~��)^\Oԥ%X�O�V�&����S�W�2��+�no��%�y�G�`�d�^�[��u��e�ݙxu�Z�����B�f(�M{��/糐��VAo���:�b,��:䧏�b"�m���І%y���'�1��E"� �Ø�k���������4�Q�սp�,m�����+�!7?k����ς6}ވ�x��7bQDʠ~�տ���ş��Z�"d� 3VN��y��=v@�&��T��&��~Y�惗��?:I�âs�HHQ��9�G��E�r`�h�'<�=K��{�Se�#����<B�H�"����]�o �<{�ߊ�����ņ�}�ܓ�*�B �Ц�!��Cq�$^�G<!k���g�G���պ��6O6<�����T��u��l�ؼw�QW3܃�5�F�w+���&�i���@W���w-Q\���!�M&�2�?��2����n>�4Z�0t��H�&�:�;�:q��B�#s�� �?m=A��L��󇔿�8�2���:��9�ζ	Jg���0������~��*\��M8��|��"��Ê: �� �.�w�a���Ȕ�����ǀal&�*�!9d��8�L�s�%��1���M��P	\�T��~���-@�汛6lIO;a��?���ļ��K9md�$��uv����������sg�k���4�;<)|54�Z�>I;I0S���#�s�D`��=�9��C�LI���p������OtF�X���8�q8<���r�O���G���d�xd���Hʏ�s�y������ر&�]�0W+~3�1�5�&.���v{,�5r��E���C����P)^�TՇ+�3ՈwE��E�!MB�oЮD@щ{����s����ɚ�-ʾ�Igg��|�	P�ϸg�Q�QIY2��+^w�'�W��#>�IT?6�%����=�]j�c���1õ����7,�ܚ���M-�$��{�P�%�y4���$�M(� }SҐ[����}�Ic��SZܢ��6�I����T��Ʈ�{n� ��Q�<��j��;p����s�>�gy���9s�^f��sS��U�F�K]zP��n�ll�u*�>~3�� �L�;�C�&��2-���P��:l��R����a�2b�C�F��	��0*�������\	K���`����z�������� ��9�V�Pa�J���K��ϗ�Lo�Z�ߜ#m��0x�h�Bpv	V�^�z�Ex�*ɰN;�^a��?�K^Wj�b�'�T<��Ǔ�c~&r^�S�� xB
����d��	n��_K%�|� x9��GT�{oB�
ɧi05�+`�fߖZX�)��W��3�D���i�/\�{-��Ĵ����r�s��I"5:K����9/F"���n�O>����YYb���5�}1+�/�"i�O=������߸h́wô�BC/���f�3��m�۱�<���
%��7dkɾ��������R8�Bj,%��a�/|��E�w{�C��;+"3�p	)G/�\���r���+(rraC��8�a=y�+�~l�D����"��,,q��y�x#���h�"�Ζz�����p3b����5��-�[f�pL��0�t�f�f	)�>ư����*�n�̻��j-���'�2�ߎ����-Mv���Q�W�ؾ������h1��ô�z�_>N�V�*��3�����Դk��������_8�Ve�oy��&N�j}�$X�T<�$p�G�j�>ppTGz��~�m�q\����L�vEк4�m���������>��mf���dث��imn���D��z۲�a��w���ˈ�����%�K��.n3A!��*vq���-��3��n�Dz����u�lW�糦��\�4�:����惖/����c�B���h9�;���e�H�CW)I���cY���΂��p�N)����z�M���x�*��B�o��&/D0}���跶��t=�	�gP��J@e�K	�6[��n�'���]� Y�F�*Kz.�d�:M�Z_S$�B�'�(�J����uf��q���9�J��>F��M>�N ��Q����-㌪B�J��['eˉ��ub���/�Jf$Wd���!��:��{�Z����r�2��^��Q�=X5���.�!e�?XS9��^W&m�q��9��K㦕��L�-|SqusU�6=��ѽ� ���o?�Q�]/��3�h���D}ha����������~׸(Q��y�5�po�&���K���ru����;Q���qj��<Q}w3�L�bf��}��jX��Gg�=r~x���5�ٱ�b��)1n�w8���V�jX��ܽ.4ْ��i�����0vy�+J�/��J�,���"�eK���p���kY�b�Y}���X���OpL��/�d� Kg�fS雸�l����r��~6"�.6�C*�1uFA7/AN�u%*�#�Msx�-R6I��ۙT�hW.j�I�2G�/�����*��8�������os������u9���&�4%����KߦQN*ʇ�՗;��>���30%0 eAG���Ʈ���y��wi��^�D�r߶)�ձ{r����y�wT"���%N��]@��ع9^���ѩq����|� ;H!��Bo�]��� ,n9�Ŀ��)�p��Z@�ڑ�;O���P���70g�%׮l��?��|\�Pz���P��W����p��}�R�;l���=%�c����9@f��F��h)Lë��_���瓢*֒��:�B�#�
��v��i�Cl�7, �T,��p�׃	T�W ~�wj4Dr6ea3�����jk��pKs�x����3���P�<re墲/�U��V8NK} �-(c����.�vy�ڌ��H�zsw;6����1�W&��3��U��h<�$}�ѮP������#a�4  x���k�{�U@�Qdt�ތ^w���i���Q�y)�r�����N���ۛ��M�s@(w��'�jT�C�$h7��f��~ύ����5�V�IMg�H�e�)���!�,�3��Jw�DS1�"Ա��(Ȣ�@��܎��*��Ma1�)5H�yz�D�.w�& �Q��D�ꚻ�efy�h����@�Y�+�u�*g:�i3�'@��S���E�W��<�u� �=)ˣt�Ak�� `�����aF��2� ̋!^�����^S��O]˄�;��z���sM?p��.�٠|�c�e�\u �%�V<���D������6�ni�.���V6i>ۓ�A���oBOn	��\�nʩH�[��ڷ)�wvƧ["�s�GK�-�ٔ�"���p�2G9��\�N��[U1���k�0�Sǈ�{;�3���S�'��W_���ݭ��Q#m�@XC�˸�;����ME�XN&i����1ɾɳY��zF�!Z�<`2D����s�f��gg7�K&�t��4k_3�m^c>�G���6�R x��Oˀr��n����D/޵/��ö�x {^E�P4����u�6N���	2F�6��0��n���2�S�:P��״�{7�\}�v[OUzO��%���� ��ن�Hg������[���9Gc��k�)i���u"�VAra�؂���B�a3��,�/�ؒ�<G���/{�?>��k�}����2�o�c� ���V�
� �2N��ھcJ(���|�n���b�:d���T�w��K5r�;�`���pMUzBz�{'�nC�2��T�N�3������څ����ق��d�h��,��a�R�q����ݹ�q!�n��܏�ӛ����-����M�������D�m��=��/��d����֛:�#1������V}���F�'|���*���^��� ���8:.�Os\"%����~����_] �ɐ�`����F���t��Sf�[�$�>w�<Ӝ3��e�q����<��1�TG1,�����Y!8����7�!9�Пl-.��(�d�	�7Y�g���j����%0���V��b���������}kda��o����.�v:/77�E�_�3Qwt)�e#�E���RW�s(.Y��c��F\�b$�9�n��/��8{&yg����8c��n�������d��U�������`FJ�d�l�1{�k��8���U,^PXKY��6�׈kkg��p�{���	�~�Ζ��Ӵ�j�r��,�v͐��<��s�p1X+����z��o�G�'
��v,���ECr7L���Ӭ3�k��_�����:>rƫ�P��)/"������`�3V8��C�mo2����a��LT��:m�TI��J�������AVǝ�ʛF
%��}�~��$q���v�?�`��fsE��U��fMF��}�[�3?�H�J�G ��_�����R�YE�(����7��!��b�m�}̥FZ^�Z������x��)~l~'�1���~��3E�F�Qɥ�4����n�cY�!N��B��wU[��Vg���悁[��Au�L!:g.&�ӝ)�_P��$�.Bb� >Kqg=����e����"��F����O���;�V�c�F:��k}���'��:���}d�XJ�i0���D�Q�ћO�R��v�[��W��D~X:�`kȯՅ'5�������Y3��
O�5��QU�;�����Pd��
T�f̐�ι�ŋ�׺Ͱ_k�����ϻ1�V��?�2,iK���%j�Tu�y���^��n�:r.�{��lZBjW��������D�P~�,>f²��@����-�-t�I6՞��4i���h�e�ۈ$�pI�<�]��߳p��!��6�pK3ͤT7� Y��	t������S��<ш����ݝ�5]}�3wn$�W
!�������0N��� �z�T��i�/ݾg&x�R�+IP�)Y�x���c�q�����7����r$�������|-���UM<M�d�����6!� �.;(+�J�'�8��r��ԓ|A�d������/��v��h�㏊������5�HGo~�G;��!�'iŨ*�cTQzz�6ϫ����@����B��s�5�Lʫi��r��;���/��%���?s99U�&=W�J�P����Ni���A�������S��Z�N&���+����@��-���S��
�?߅���%�%��k���g���`-|;W�:bz���)i�[��Q�%n��P ټs$��U��G�g�A���b�ӸN��;Ae$�O���T�X�R�pk�j%v���b��9�/���0��~%隌�����`��d�z���d�9fkw="E�Ů�Pk��FX��ǈ�5��Ws��=���Q8(H�7�_/6�&YQ6�3�כ��FQc���~�/g�v�8K�J��C�̋'��[W�[?�~˯���ʯ\��k��n�}sjrYwZv�7caa�0���7e\XQ��9_�TYC�$1����ﺭ�����e���}^h���cm*<AJJ��e��Ӽ�{~Gh@�E����:L���z�5z<Yx[D�����i����Y��rfj܂`6u�
�R�Wǩ�f>����Ͽ��3Ϛ���j=����|^��1��.���]�*���q�R�y��c��F�x(���Z��_g	d������I�zI�n'��4!O�����������ܚ���5�.[�m��(�^�z�+�MV��[_:�ܨ�8�_j*�F�dk�_�5�}x껟)`=�S�3 �t�5���c�T��{�a��vvb<��ɵ�W�:e\�X����x���[�qg��D���+����|QBÂD\\|`pP�~ULZ��wbbO��!`{fee��CoW �V���3rСbQ������fŊ�������X�~Mt�bQ�<�zP���C-Z�l6[K�,�\&�k�a��RR%�SH�eJ���������JH�Q]��"�A{	���G~U�����3+'���8U�3�?���K���1�@�]��Y�C�����1Q��,�:�"X�8z��ΡO���Z�,{�l���-4տ�H*��P$�/�۱,��y�j�S.%��ͬ�ío����f�1�We��'GWqK[S�/�]��"�k 9[�P���5�s}m�p��u�	3��zMϖ�k�y(�K��� ��`��Q`J����~q��Qd�VW9�/�f�-˥d�/^��x>�M�K�ݫ�s8�zM�P{O=@�	n����8i�Ԃ�;pw�V��%�F_�U��
��>l���vNf���L`�:�3Ш�q�Φz����م�[/���ҟҧ9����H���iIM�3�%���h�}� H��YUH+c&'��)Z��~��-f�׈#֦�	�ZOYKf��s/��:V�Bs'ɹnMsR|�&��#��s�7�|YAe�pG���¼���
z�&�«F����Lᡈp�2h�녵�8
���w+*�KVC���-}�JO�n�E�IM7�8�Yd���A8 ���evXɣ��c0�#t@��;.��w�ɢ�HO��an,k������P��-�EC�F�><�QcU	���^�ͬ&Q�3`W9"����k�r���!���1����d����V(�3����խ��)�vR�QF�q�k����x��5����g�`�ԁ���5.i�3?k�'��?�������c����x�,���=7e�8w��P(T_΀9L�KKANb�+�h@g��?<:��Js_�s�S0���C��ϳ��~��Cn�xh*�P;JJ!�0��އ�g���Q�� ��Ktd[��4���Wd4���2�b��YYS�?���4�{������=���?�c�J�t��� cK+�B+�I�6l��a��i'S�]��]���k�p5���zlP�̥��_8�c�ڗ�4y�y�<�d�z
�*�k����lϛ�S|�x�g{��X�J�TZ�eej����=jQ��%��*�G�+v����9���ef�������a�fS��<���џČ�wػ_QOWnPe�o�Y�ƕ�[�,/ۀ�<��Ixx���Ɂ���e��t=!9�f\�8+Ѝ������.n�Ð$6�E���E{�,yʆU+B~��P*��HW��'��zG��(ܝ�,�ew���mg���k��|~� �&8�Ey W�80��e���ٯ����S�9��!-���t���)�ծ�6��aj�l}��@�>���QKW__5:XG����>�*�2+;��}W����i�r[)z8��Y�X�|��5����RK�G�H��F�2�����,2�Ng�Gq�J��fn����l_�p�E�-�7��sR�o�i�h.���,���HDy��,��S�� �u��2R0�.�&���w����dh{��9�٣N����c�����C�V��C�-̜�O��	up�/G��E�Sl�3�r�D�~���+&����[T$I,���y����w�k��_��=1{�|�����U��46�>��AFM����I�o6-=t�x�y�w���W*��-.)��؂{��t��e�G�Э��Q�nA&��/�E�R����m������Z�<�nT(-�r���Jt��q�Q�L&���( TXçA����{o�(����:�;�C�|�~� ���xb�H�]w� ڑ�o嵠X����ȭ"[\"�m�N���`���h$�9�_j�1���56`4�`���$��#����3���TQ��裎����G�"�Lf�Rͧh�5O��u�-*�*�� e�������f|�i���Z�B#���T���i�Z��O�j�#�q���X��w��Y.�>�2��<W�:���t����kKBѻ8���D��;�(�ެ�:��ф$��H�σLx�/� |g�{i򈨅��|���>2����z�I
|&����s��6�����w��3��f�E�9�?�|i�G�m{��F��q@��c�~X Iqr�%�m�[)�!=䙂��u}�8��Qs3O��EԤbf�m��5u�}2���'E�FJZ��ѷ�]մ��d��4��H5���z+��{9��X ��W(t����z���7��h�/�-��A��u�郕T���
�yP�hΗ`��9�؝4���D��5�̜t/9J�M�L�m�?!�*�A���yw������~�������Yi�losvD�F��0肉��%Ŧ���d��J�6db���3:p=��{3CV���"�{I�bs|qpCׄ������E��U��^@���3����<����!���]�Г�ϧ����5rX��c�8K� 2v�Ywb|d��Q>���騇4"%�r�0òبK��v̯o���k�\r�}�H�?��;�
>8�ª�v�M���$86��o|���57t����G��ٶ�}�T���Y�6��*�����L�b7:<?��ɻ�>`����{f��q���M���u����~��O�qf��>��Qk��V��m�͸=!��#��}�F%��r��>**��򢦪����&_�i����c����t'�1&�.ȍ���؇6/�V�[��ߩ��ě���?͉D��ZQKTW�w��]�����Y�1�G.yuV������8��ݙ�eQ��Zv1��r#Ew�}C�.VC�ma*�͜��otp�+��S{�oo�;p��,�(P����A�š��=��6'Iѡ�.僧nowL�r�*��!�>�RkI{{9@(zV�F�L'�$�J����{�߰��ac��^us����jij7�57���<w��统L�R����c}i����7��*>����26��vGN������*j-o�=˵�F7甤��Zo[�Ƌe��Ug�,V�Ͻ>�i(i��).���m������:-Uu|.9^//�)NqqKK-��.߽n/P-������@�^Jͅ�آ�v\o�Rl�ˠ#i[g��ʞ��G���Xvo"��o_�v�[{eo��dI�[��edTMr�����=�8��B�on�p�$����+[?��"i��K3$3�o�
�����S�d��2d"{�_<JN����iG���
1�-�抦�;c���PH�d��P��VW��lvWū�u������~�~���>6P+�^����)&���^�@/����&{zǚ���`�-���axa����+6�#{{����y�!֣��1ϒ��CS_r�������=kN1@�>���C
Y�D�SQd���N��������� =*��� �y�A�� ��ym���������g�Mm-�L���=<M:��,:���:�U@���E��_��2Z|7�2$���}�� ]�iȌGsy?��iw���5d�m��Z�i�@��珪���n�z"�#]z��_�mǪ�S@�+ ה7�)m��.���Xߛ*��j�q�x��9HMն�=,>h�������B��6�\ݕ�IoпcI�A�x�FZ���Y�D��s3�ua	=� ��������)@�0�j2ӧ�[��Wo�L�GL7F�x�X"o�F���xȳ$�Ƹ�3`��-�F1����+F�͉�K�t
&L��.�� y�l���Y�k*��v]�%s�W����rv�ҎFv�tn	�(Eᤙ4'�Q�c��4���T�9��/�@�D�x�R/_.1�cmU˹�߃|x|�|�X{�嵮R�ݿ�E
�K����	��
�V�w0���^ނ���k��&ۑyC,�^�C����iF��0C6��:M��TZ�z;/!#T;�tt�\�c���/HŻ��ZL~F	�����v�z�|����u֤Ư���\�
�ce`��+�>D����W�ɽӔ��	�v�g|+�������d�-i]��N����D�e�Xm�Iħ�F�[}r͹j��+B��^����zF_�+ɫ�xp|�(�ߣ�g�3�Maa��!x���ª��P]7���`���������T3�'*���|=e+�4�56����K�&ذ�MF?�5���:+�����[oI|��r��zdRy�p���aX��:��y)��o.��C����:��Eɦ�����͇�`]G"@��r���ֆ���Jz�W���5ߜ�I.��۠	��_o��Tt�h���)˃�}�;�����ǳ|��eȄ�-���y�:E'���-i$�Aѿ^I����%��H��������G�!~+/�f���;��qA� ��`/!ALdGs;ʾ��d�ߏqz$��ȼ/PLe�k�kKf=;B�}V�
�[���l{-��	k("��z.qz,�Òk�8�#��\�՚�b0*ry1G��9A�`���sO�h�>���}�/�F����Nf��ޛ _	2�5��I�"����;�K��-���Bp,���*���%eg���1��?�;Z��(���)(N��"3 �{Ǔ�����%�iV�Y��?ͭs\={�\.�V�B��+2^6LX��
��u����>_Q��Lw`,t��c�H*�;{-��Y)d�)��湼1԰���A�M�[�+��Iv~/��M�g���)c������,z�dH
��%�Er}��zN��_4�2h�}�ʺ��~x��f$��1H�,`�r�ñ�ޅ2aȯ�?j��yhK�:z�H���:��-*�ægL���:;�"��H�m���J���ֆT�&R�w^*T� �i�Ղ�ha%QԚ� ��e� V������a��H��I��r��[�}��Eb~�+�e��zS�-�(A�<.��1� �$b��j�3忮��s���bn���GB���+Ө}<�g�N<��0w�Y7��H/��Xš�KF�k�L�d�573K�Y������U�!h/z�[�p}N@K�sQ�o�3r��pJr�U�wɣk��ڋ�!.���xp
FF����v4��;��F2�v�Ӣ�EW�����]i���:+�u�s�Le'���������A�n�
p���7j�ՔF��(+�.����� t���PEk�RN����}��7���Y���c���^�_@������G{�� �(�+���4�.>���]�t���s;�h������6�����j��Y�E�M�qLt�6�4#�m��-�٭J�_����}Ƽ������Ҁ� ��}��)�U\oKQfm�A:�IA����^��kD�}�2 ž�����qEx��K�ٰ��&K�	q��~��꼋�vNH�z��<Է��Y�"��=ˬ�g���m^j���:�Ugj�g��/�����i��e��+T��-��n'�1�:Y��L1r���#��:B����S�\V��ӇIkE릶�V��`��p�gp��մ�1�lwLYә�6����3a�P������m�^�k�'Kc�Á��LluUi��m�@u�}�𞁎P����-+��l���i�_����AAcZ�n�a�3�k��񖷿d���ǅ]�+�'�Gm�_�V��(q
�4p��],L�؞�1�dui�Y���^�d��������l���sE}���o�1XtQ�����~�����m��k�ӵ3j�Ts��Gl���� ߱�5ѳy->?�iG �N������>��G}�-ec��il�����t^iţ��c��PfV�����z�U����AȽa��(��Kعg�r��~�X�����̔���s3�����1�4�LMQ3G"�9��"v3�[�I��r{�nV�M�[���8��w��~��Org<��$��[�$ ͹hk�I�A`�hk���;N�ˊ�(�h7�P��:�.c7�fCD�2T6�L��s{}m�#�ڙЫ�[K��:�-��.������.Ẃ.}�u.��	%yǃ�̬P��1�_zWi��$[��C��^+t���
�y��f�r���+����,��%�jbr�����xx�vK��`��D ��mP�o��CJq�,f�7�P�z(�QeKFܫ�~�$����"E�bZ�gCW:�q�*C��$��S�����<����}Ƀ�l�0���9��o��b;F����N� ~t�
H�AS���bJM�x���2, ��%[͢�,�=�݄v�Lem<}�{�1����Qf[��Ԃ��$6/5T�.鯭e�R����0u��<��	١\�%��`�Ĵ�0it<V���#�x�G���7k��e䄍�U�;��rѦ��:��:k3�'_+Q���Ӷl����{���*#��6	�y��+(������6+�K�y�@�3�.�:�)�{vq{�ʋ�4L���Z�t{x6�f���,Wf���h��T��fj0���I\�]-�� �8�u���>zd��,��<733�t�q����8C/�V��t��|����a�<�$2�j���ȅ�7.������zDR�YP���7����v»�nO�c�F�|2˭+מ�_�oj  ��h�^j뇸4��ܸ	��e���Ʋfd�B�m	"��t�ࣱ@G�
�0�����tL��*[
�F��~���
cv�W#�=Pc@�F1����ǁ��brr��PW�v���Ċ
;P�UU�+*h��n%B��j�	9:2�B��43��-*
>M�]�Е��:�!�c�y,�:��@�5;N%�cl�?^W�gB������STZSUN�E�6��/.),{{��Q���]�������ހv����5BF�깵j�zC�ޱ6��z�3�;�E��ݭ? �W%C��wM�W�k,��qc�� �Mw���*-/�P�Uw|�޲�!di^&a��F\�ɥn�B�E����w.)���n�3�qN�-���qG��H ���^eA�.��������f�Aj��1��:��N}sЊ��"�켚���a�Ɔ�X�-��������4n{�-7�R**V ���B����ك�Ʋ�mR��vW�=��������tmj�ݼ4>����Sd������!'T縖-st��$��铓!�N�<M���b����3��&�eo�;��c�ľJ<��F�d<-#;�^�H�k�)X�ܡٚ:�]�v��@��}���ƕ�lwoj�M�J�W�V�P��S��+�����#�-��
~:�!��Ԧ�8�<����ͣ�]�}?��3��*VE7��\��Hj����Ŕr�J�4�b.�y'h���W�*���?����:�����3Q XҀ�)��Y��";Lv z�ث�;�6^�j7:�3���N^d��`U����s���N��|=3{��6��`�qPV���r'�#�ʼ�P�U��LUɀq��������5U�eo�����16��ܱ�X�=�XJ�������|;*D7�&@.����Y̲� K����?�lt��M:�4�x=P��\����l�4y�ϱ3z��3���'f=�:U��-e�q�M[��F����03�����ָ��.L����j�;�`Ԣ� ;�����ߠ�[&��H��ر�F��DjO��Z�u9ءZn���MG~��1�n�VPS����Rh ��t\Q��Qw��`�K�ٷ�����|a�
n�d�v;��h\w�hC\/:݈u�5�M�%R�x��2j�yA�l�e��L�4�N�8�hq����xD���fTO����_ٹ<�骥����,\SZ����V*�ڝd�{Z�����N��B�+�ö.�����w7��a�vt:1��/t=<���|S���������6TM����|+ѹ�ͼ��ſ"����m�צ���EYW�>,u�ʮ��Me����m�
��]�{(<�o�ƛ�|��o�O����P��g.;e.�(ʐ;=.�-�s�'�:y]��QO3��eY��t5�2�:�Q�CC;."�;P�	a��� ��Zѹ%�� x�ʻt�Y�{ƣo��)���;�V�5榜�ָh�l��up�0�LBcݔ.�����}N޿�+_�����V�׊�%�\�δzW\:�'�B��pcp:������(���_%�(�x5n:�闶m�T�lFvi�A�K��KoA����[;�*2s�N��U�N]0�ͯg8�1�޼���L�E�����/ze��L/.�3Z���j#���o�����H�mv[�쿸툺3���S�5��}Q��
q�J�F6�T�Xm�uO�ɠ5r_�H�c���<x᷒�����Hﮃ��G�W���E}7�=2҆��H���t��ʟ*OO�Z��r�����w�(4�.���D�/�뾌�����<OK2<x�cO�Q�~�E��U����6�43sPԶ$�br,'.�)[n��"uzzx���h�\,m���AGIcv)m/��j�u��ۮ_�l�Т�tձ^*�<mS�Q�ϧEy_m�k����b)^�Vf�M�sM�AP�Ͷ9�r����7? ��[U�-��c��?0��C���>����|��s�|uF�W�.�5��t�ÊJنgo03�@)�P=�
��ԕK�.a��r.`�|.ǈo\��ٰ�)��:�il�y�=:;���V��Y���o������$W�H|������Sr����;�$��ٷj��IXXP�ЧD���ޖ@�K�l̬���xPS�b
�3��:uk����C�q�5�� �K�M����f7pyW���+�kf>��ݸa닗\��/y�,G��/<����\=��p�yv_�����~�-�ܝB�{(U�25�q��G�!f�9������1�1���}i�k#�7BȦ�h�����Be~ �Y]����:���P7�$0)�kxH8������-`�ݢƗ��2�
m	�çUq�u�;6�y쓵ֳ�d�F L�_�^v���5ͷ�Z���`͞����Ļ��պپ�yY�ar �x	q���H*Fb}*�I�J��-�� �6u�w=XsC�ve�Ӏ�q"S2���\���_=�{����Z��2��e��*d�/F��* ���W������ƈ��lo�ۛ��*~��,p����,��]����:�-C�8}Ϋ)߁��3
�� [�����%�������3��&����VX[d����Wed��s����ܓ$R�>��*���v���f^�U��q7k��Y���>�������.>���W��W�M��q����Y�t�a�Co)
={�y8n�OGobfo_ю��5/��!U�N,$5(�W�a���n�x
�?^����Y���uI)��d��F�sX��y�͌���OY���L��X��Qp綿����_�E���^-fpIL�����|�]?t��:֫�������)�v+�N�͟7�#J��Ǫ���d�溛��V��o�J�g.g��!���m��7��
ҏ�zb;^���΍s�j8IL�W�6}/��L�A���GN�2���W9�~�[���΄+*�?ǯ�'\ҕw�u�K�n&���4-0�;��)L��r���]�#�G���888iȄ�+�3v�j�?��:(��EO�@ @	$��!�����������wwwv�������ޯ��?�z�������>���+��6�I�̣��l���g� d4���08����)�YZ��@6-x�|�<�N�o>�99��(X��.����F�)73�G�K5Qa7\��c�D�P!%���{�� 1Rk=� ����
ޡ��ti�u�8v{���.�W�Ϋ�fzIyS�+�_A�>���C�����s^j�w�ٮB���u�$���*$S���-��8�}��������}�"�-�Nf���Gv���)6�ཀ��;(N�Q�k��M>�[6]�ߵ�3]�{#\�����(��8�ɒ��P�H��w�6A��5w���1�^�ci���Tj����}k(�\c���,���J�t"��-�� ޒ"�<�$�.�e�7M6��(f�i��"]�c|���[詘��b5��W0N�2�Q4��vة���~�*AY�(���wO~ߗ����j���)z�-`&�7�+��`�9mW���0��Ԍꬤ�棄#��TR���3��D�}"��	�gF�5���ry~��>;��e���/6��'�=ᛆ��MB�.�2���ȿN[I,�Դ2�	�����F'蔻��<j���W�nͿ��n�E��q��)_e��T�h�ط�{^Ё�J��Sy4�;~�s��B��^���mlx5G��,��k�z�1��o�~'U��O­w�s2|����aҗ���D����橝'�Ț�:(����ٶ�}�OR�Ϥ���v�ڇ�Ⱦ<�kZ�qVG��8p͙&�Z�T1¢K��&��'�=���wE7���o�Ԧ�bb�R�I�!Av]L�9y�e'�H��xS<���*�:�	<$�~M����"ob �k5�UGp:�fh�Ub(��a-qv �Uj����p♰I�r/uμe��O|ĥn����؇o>�-(�~�(��o��P�M��`��z�C�UYwSr5�(�5{�yj�r� εI�Ո��Ҝ!{O�we�1�9�����~]#�a���:MѠI��hmZ^x�T����3i��s���b,�tAПV^��b�+
�[x�O�m� ��Q�[��{�},T�9��:�tp��R�^��F��/.��jMD�cy�DA�I�B��m�Md
������٩��Ax�����>BQ�ޫN)%˅�s�C��xe۵�b���{�(��o1��ck��omD8.	���2!�&gg��B�����,���d���4̈�W��X��B����t5�oWT�9���������Ȣ���K?�[��'��߆i��(_�x�k�/0���=�:(�O��ʣV
�P���S�^��Y������]&yJ�xgK���o�����w��"&��rW���٦o|S�ً{�-���-yg[����F����z�`*/�{�u��ɳ�q�>���O��*��+H���W>�ŭ^9DL��;[O���6�s���k�G6�Oy�1	o�Y���--�(��	�<�@�c����z(I_���%/v����/��h\๘й$�W}�]�ܴ����p�dfue�w���Рӹ��;d��c���M��l���#
��{�Y�6�H��<�(�M`
.�$H�J"ptJ��<w<���h�n�)۟%Vh����8���I[ +|y�0��w�e:=J�|zU�*�޶�5s��K�Fn!���XK�m�5k�"��b_���3#��*a`��d�!xq������/�m�{k*��L@�:�gXf����U���.�Zi�������qm%e���;��%���G$E��[M����:4���*��Zg����|]�����4���ʼ�u������L;'e�3@���(ֺE��Q��QW�Pּ3��>rޖi�m�@������bF?1M2�����X�P�$J6I����^k�,����9�%���(�M!��V�a����h����y�M_�ʝ��A��l�K�H�a���uCy�5sH~���9c�w��肾������{P�0��\��jg�gv�؜<~�^�HY>4���eR���E�\	�#�G��M���E�22�kK����Ca���U-�Wz2usy�9�c�)F�uވB��8A�!��+����nKɶ<�ǁ�6ĵ���B�)8�PX�,be����O�e��5;�.ZZ��K�Rw'����Pռ�"�NxtU�25���Z��LW|r+`�ꚼe}H8�r��v���#Q�>�E�d��>~-̡D62L�<̖`��RKc�p���ӫ���4b��xش�'���X3L����<�~�믽v�0��~b1�þx/��Uh�$H�i
Ҽ��ؖZ�6�W�k�k;
y̛�dWc�$����O��(z�2������ S¼ ������K�p�:Xm�]��4�����#�l��N�un#�c8��skw�>5�w]�xo��3�V�b��������#o���և�.�M�u� 03=K&�wS��Zbp�JRq��y���6�1��C��ϱ}_~�,�dTR�W�0<8��(ʹ�Z0J�E�OQF���	��4^����͊���%p��x=����e4@���onpRikP@JG@eJk�� ���ȏ4�3=�+��:���e����~&�X=�r��.�/���f��(?O~���@6��R��ޡp�7��Fr;�Q��m�NV��$�|[��]cY�S$�t�`�=��/�/� (	���U��|a���j�cZ����
o��,�����hYS̔�x�e�
�Ԧ�wk<r���-�cT�Hg@���^+[��6!�߸p,d���x�Q-QK�2X?�(��#  6ؖ<�pE��z��V�*J��UK���r�܀S��?�0q����b��~2��YK��ZGci?��r?$�Q8�{�za�}�l0���uN��<K~��ϔ[1
$[^Jf��h�k{�eE|���nw�Tp���w=7�9|��%�__A�M�u�<ǉ+ke�u���3_��hG��	]��V�y���x�m����oU��)p����0��vf�� �V��ޛ�M�:����G�zG���]|^��|&��.�/Z;�[�tk�f�0�����d��*Z@�/Ï*'����ne۽5�-U;�ԅH�ѳ[�!s���P��l��"��)Z�UCV��F5��P8���P��,]o�X�Ӹ*P�����(1����ZÛn���K�nRX7��k:4x�Fb�+�r}m2�+�;`A���\a�����Y�Ϛ�Ӳ�X.�8a��;�U�ոV��������#n'�����M�ε]��rԄ��j�֛;O��$�G�?�7.�h�=�} ��*oz|���Ǉ�eM.�*�5ɯn��+'��gQ��*��bk\�:���L���]�>�:N�z�.�0�DM�V^<6�n�=xHAؖ�ˬ���w�xQ�Ƴ�0k9����^C���bo���Uk-ooa��;������k;�B��5���7��3&o��Sۚ�a2�ҷV�;�9��k�X�ŏa�C�mK��_���)�:��|Ο9)�	p�h �;	����o~B��Է��'�,C��o�`c�-m/�N[����]�ak��<�%謊�(���ڐ?����A��B��S
��GeW8�9�O������]����U��W>�:�!4+�\{�klb	u���J<�Dd���uߦ�N8�Z��*C}��n�N��|v"5�؝��O �ϤU�hg�S�w��Ii���/x��E: %�;�:hr���h���g��[k��oI�"2��?�����lp�x(+ޖ�86�]!��Mk�p:됸�oD���Җ7Ȅ��~�TRy�na�|�r~��-��Z� K�|| x�ںF=�ɳ!-���`�R`�8�l����b'|�'��y�"��3�D�
Ω�Y>H�$��j�2��P
H��^��I%Ԑ��S
s �ǌ}��!=�\%�P0��'�&����e�/�3Њ㗠_�(�,.�s���ꛊd2qb�$m�� _MFG��P�\7�M�'s��d�}�Mc��ҹhH�͕a����c���#��4�KZ�rv ׾M���
�z�"�/	~L	�22VU����Y6�qc��^��r}ֱ[j������er��H�JO<cʷ��j !3�pj*ĸ���(l,]h����Ր�D>&�ɲ�MDy����ؔ9`9���P2���u
�~+0ox��+Q������t,��S1�/ٕ��2��p0��,���j�_��8���aY{t5)i-&~�5Q:,	8Ī]S�O��lϷ��qA�w��&'�"cd���}/��5���ݍ��������VJ�C!g{ I4�3_1�艳���-��珞~e�5O��{��Kfv�idhB���V����1���ݰ�c����B�C����٨�kX�6¿@����9��7P1-n�A.�k��'�o��V�IV��C��OA����<3�ϯe�����?�~�y!��Rř��M��(���y�����k��_��>�n�����,�.F��0<V��f���=cv�e�׫h�߹H��!#˔�����kQh�<�A��۞՟�%Xa���I�;�No��?!����=C��ֿN">:��-��&U���&t���m���'"�a��s���NG�K��r2s�<Iګ��ffy/�_*��n��o=~�o�2�~^/��\�E���3��=���5���%��*L%ʅ&���)�R�l���ч���@#�]@�c������Al�I�Et̚��!�;S���D�~郥�6��Ǐ�,]"y�y]n���u�cY�\K�P��U���{�z\QH�?2�Z7E�r���Q��Ǿg�����s�e�Y���NG2�VN	chg噊�E�3�$���/�����S�[R�A����Z�����%��ڼ>&���GdS�s6ng����c,�+j�n��q�lH_��x����&����h_%U��yq+@��B��r[0�c&��~�s��g�ᘲ�g�#��VL���������~� ���	ojq���4��P=���%�6��G.�8����CЗ�$W�������G�ʀ�(|K�|lhj%h)/T�(+l�"�O�2��V�2���+t,H-{�SģJ|�M�[��,@|�kE�������tmP�m[��놛Q#�/���^״�c��zZ1��b�z��}��s`�G?oĊ�.�R�d�%>�/�9
�Vy�5ї���m��:&���Q}%��z�w��ڦ{��J���f�?S|$C�ZYd���.}	S���'"�Y �M���s�?q��.fa�1�U[����ס0A��
����'��D(Rl�k�3M��_��훉����v�d���_}��r����?:Կ���n-�ū�	�QS��ƕw��f���b�ab������Dy3���l'>Z#Aآ���O͗Tp�o�:g���t׿�:��~�)19U�t�-��R���R^�<��enLWv؅���|5���];CeQ2Yo��;��.5A��gS�v��y��ER���L;rI�p�,�˝Z��wz���	q��S��G��Z3Ͳ�����������v�b�&�;1
���w|����8r]��p�v܀�̗�ԯ-��r@5ښ���[4�l�1�-�b7pE������O��ڶTx*p�jt/�m�N�gkpt g�v֘�cv-Y=ǒ"N.CҬ/a�EcSI�}�RV$Wo�n w�h-���O��ۿ���:_��r�r�s.���ep��'��wŤ�ݡh k���_g]�P�V�9��G�8�S�vϵ��T��u�l���Ż�_�?$����5�w�RB��o�=uWՊ}lp�f��D���c����q��H���hF���خ�Z�/���o���&3�-(7I��Ƃs�R^	��%��>������ۨA¥Xo��_oC�&zy�4՜������/}�ߕ��$Ic�*J=oT� �ѳˠ��}2��s�'��U3��c�wN�-#����~��Rr*�H�W����Un��ۼ~����9Nğ��o�(�:f���?�<�-,���������U���X�������37�����r1ޜ?�;���Y2��7�`�jl��UM��$m���,��@}H3��4�v�3�h�E�0!�D0ǣ�)�-���=�����
w���Z�)��j��?�@�u��4���"l�PC��d>&8�a��f�=n{t�ĝu�X��?����������Wf7�%s4����dn((�P�. ����B��t�H�f���y��0�NQ��*
}��ʮ��[`����В�f��TóU����5�"k���݋d���l�_�龖�=�֩u���Jϋ��
Dj�߁5��V� �U���2RL���|�;��}�Z-��J�A�b�|��uh�����P-�2��m�B�2���D�c6hv��m5�QWf�oX}���6;�<;�:{���f�+� ;Ev���CQC*U�;U<��+���^1f�W&[۪>���2'_�����`|��-�S;�=�NCC��@����D��������:>@�t��z�m�;8e���g��c���=����2�t����>��gV/V3��⻰���v�j�� ����&�tZ|2�6hPR��w��������j>u�L���� ��?��#�Xv�"\�N_U�:���ͽ�[o�3���MO��lګ�9�������t2�VN΋(��t�X:�lV�j(�l��4f�W������?�Ƣ`�-���o�O�|Բ�y��_��l�3����-�;-���G�D�Q�ʝC��zJOW
/I�=SFZE��"�3��F��֞x�H(g�/H�����j<I�7� ��֚���$�]�F�]SS�T�l&o{�'>�6�X� �r���Ů������0�K;�����D��3�E�"���w�0�E�s���4䫹%(�͑�6��C�b^�'#�;�K;�U��y[j��a & 
s�E�E��e_Հ���*:�>Κw��N�&*��Z���̣cR<T�����:��W�U���`�������J�6��M`�M�� 93X��za햅���,��:l)�5�f�C�ȵ��p��V!U�P�{�{Y3cgz�5k7�yȘ��k��o��0�,�ae�mm��	K$� ( ��m~?�
��`-q�� >��֗��'2��L7�_L�3��N��^Yef�o������qc�?�jϬ�~}I
c.t��G[LzlDDЌ�o��g�T������er���pK0b��7H-��(> 9�L4�G�DV���.��fwF����OD��r;�(���{Sc:��W�ڥ�����&��xT��j��-R�f������Ui(�rp5✬�����O�i�f��-��ov	>���|�fZ�,���~��c]����U����jdӔ��A��
c���h1<AI���˒.��y�.;(*`�[T��/I;�'9�o��+�v���F8'�bX�f�t���QH��~Xb*����e�j̢M64�8��N�n���kk��J�tN��⁼�G-���rW�|o��$7�-bT[�����ihpߴ���Y���l@Y;p�p�qW��e΃P�<��}� ��������!��n�K?K��{�.�N*��}e���7�=a$�K�y@ ��
�h�M����o��d�>��67d3�P�T��'���y���}����4��O��=%�f��Xք�#�U�w[��]Ɇ��|1KS*y.��O6uO�Y66S{���F��Ґ��-��$��>�y�{81)/�&��`ːщ��VJ�j\˫����ʷP9й�xF�,v��/;d=|�?�W՟����}/�Cq�]�q�6�r�%q8B�G�L�
�VO�[@5Y@��b�8R�sE$�%��nTei��/�Г���A��?=�<?�� v��,�;����{(��-\^��k�p��U]z�`xT��֦����74�R�I*v�Ӣ���p�VNG��5�������!M����)B�S,��(�ҳ���^�7A�V���U3�H����(Ҝ�-dkY������;wѰuJ��l���S�^�[�I�Rr�t��[��#%��8����%���a��p�ay��"�_c��f:�r8p�PS���f�ԏvCC�3~�a���.��uT&R��o�S���f4Zr>��f���U\V��6����)�`N��c�6��N83B��f2�o�.������*9v,l�Җ�`>/;���6߷l>FU�d����m��gMf���]������(��|}=�r��)+��P�IJ�:R85FxK�&R
�È㺿g�~��q�F�,[�_!`�J����Msu�����LPz����`��7l��f�����q��IA3k01A����5������1ʿ���e�%.��3��.f��&*%$i
yo�~�QKUE�������gI9���P�W�t�>�)��I���}>f���ٵ�좌u��}���������I���OXX �+�J
P�������|��"x��i�������4b�����
=�7��S�i3u��I�G���m�� ;�7������������-`NP���L�;���<_G{T,�����u���p��a���y��@���,�]��ۘ	��;ژ��I��s8	��ox�v��cN, ���Է/�t�pͪ���Z"�/��2 9vx:�|�#����������N.;�L�'&+9�{��K���y��j�ܷ�rfˀ�K���� ��ċV���.u�rtGf�]g2�E�e�.,'���6��޲i�Q}b�'mK5���ld��v��)�����Y=~���y�i���>q���PBbB�C=�4͊�jW�Q�)����5���ſM���B!�ę�ðj��2��&E�W���\�������j��G4L������uM���ΒZ�B���x�Ќ��W6�EG�ok�f������G|�^u���h�h-B�T�t�0q��W+�{�����ؔ���e�o���!�usƪzO
�r0Ǧ�����VA֔Τ���7�(�t�&:�)��y�o8��H���MK&�	\�<i���^+�]����jj,�mu���@�SY��'����X7ِ]��%�O��fF�["�^��1~��7�?��{�w\K��EK��_����JL&*�����+'�� &g7x	�2'��ސi�)Vv���ny�.H��G�c������̯4��o|��D�1۾Ht4��?�n (���d�LHc�X��&�%;W���k
������X0Ɏ3�E C�4ܝ�
't���C-����du����Բ#��p�w���K��p+C��;�$����%L㑢O�$9���<"�抬��Ƌ���Bqh�f�� 8��zi����:���������f3�͇[^XL����+�������/T��~j�x���=�9S�+8ĥh	��֬E%Թ�9�Օ"��r7~A1���(� O�E&,�|;6nj�o��i)Dg&�:�W�n�_͕y�/�s}�����ɔ�fvF(�4Rg}���~�w���D�o������֢�Y�'���Ϣ����D�w�B�»��V~���9����]|�܈M���c���T��\�{5ƹ�t'�,�k����ڬ��.������ׇh�!(ʼ�'�sO���g݃�G�sݎ�81�o秊�/�)<&��X��gF�7��֕��ٸG��[�|���;쎡�dT�Mv_Ha�
�_\�K���/�a�4�x1MdD=��#�8&v���G 9=Iq��pl,3�����Qxޘ�9O���m�JLZb��J��}���f�s-98!��]j� ^��*�5M�%bY�r����C�l����=߳T�]M�[���=3����U;��;:A�8Y���at*��l|+>�E�GR�1bV��}:�V�&-))�+b3#P��Z�[O�o�-�f�jՈ�/�c�~ ��q�:���3&�K��Z�g�1�҂����ć|��U`�N����`7Lf�Dq������%


}D�`U�c���Ed(����3T�k�r��Ω%��8f"���sh�wZ?^��8w�E���:}}U��e�ԣ}?����>ߘ�[N�~/�:�nn݂{hu}�SR�	�9��/�bqf�0�)[b�+�o���-��`aa��+
��1�ʯ���t���F@@H6��٥��_~�n���<�P��>�������;�8=��w;�kB�i��V�߯�<nM�ڮ7�waz��=�j�wW�d���@yM�߳��QPs�}ss�����������r�+���= A/r`hhk��P[Yˋ���f���̥�$Ӭe]�d+��iK���H( �[E�7�>�X�_���f}�a�ና^*�*��P����?�@�01�<��$�ps{�+��5�[~�NY+�0Y?R�o	/\�#�aB�
1lҚ����&����:(ͭ�J�o�������$�8�;�����v�iTȓ$*�E�\���؋������J��WY�b>t�5�6n?/���sk�@Ǎ�4�Vዊ���Yf�����`���M������y��\��HɃ�ۤ�՞���4�)���M[	�$�)�?��������m��>Wz��	�����͆����u��ݨ���DԒ��g�ffz��K뷰蚮�D0H~�9��<�l���g��8��'Gy�h�ڈ!��1"F.J��2�����r����?�z3��;�l|�P��l���9/��s�:�����UƘ�Z��M/�ž����8�~�VO��w�3�{�q�ɞX���ƣWx�a+)�c�ϓ)%?{�?������uX�-$g�ڈ<�XH�����R�JF�p�] �ۋ>jp_.U9�vA0O��m�<�Sq��y�hDm|����I�'��4�m%�۟n46"ɰ�V�N �#�ro�C��l�H�*��P>��y��!`�����{�e�2%��M&bmE�}}t�ijnK�2���N�Gӿ����dT�j�[T�������+^��|����<5X;e$���.p�s/�j���՝�}%�$��B�9���/RR�L1�=�<����^yբ��p}>E�#�wr�arS��|�"�8�(����+�9�$���s�,,����'��R�P��N!y6��9���}1ι1|��<*��%H\��~���#r+3���xx{\	��y�}u��������9�T��^g�ÊOȐ�RD��������`�~Ԝ�b+��_��2��ЇY{��,��hU�W�nlk�TM�k���c9�w�75���\��YvW�G�+,��j�-�[�^��|�uK���9��d���S��bsl;GC�H~��-`����MZ)�n	��!�=�F�҅�͊�-w#:�[���b6-x΅nH�p��Do �Ĩ���jĪ���O
jƸ�`J�Z��74F1�)*,�6��>|s}k�6p��:��YY�&@L)$C�0��� �Z�^z]Ҿ;@�ʬnX�����{R޻�����hGb-D�slY<�eR�����V�#�Rr�m<�`Է� P��E-�,;^ƅ%`��R���e�6"����g1�ƽ���~���7"��TK�@��"�t.fla�e���U���Km�E��p���(d�ۋ\���~6b�"��'���P�����R�I�əT���2g0�('c���k��q�$��ٝ�6��o�b�l6پM���Mk~����^����pm��8 ��$�<�W�x���<>��Ƨ��������"F�|s�]�F�����h�q�m��C,]<|�NVkk�Ƅ�I�qfzq5��v�����Y��z�+i��Ǥ���-vԻi�.Ƅ2-�o�ud��,�Y�P	���dQ������c���	��\|���T�4�rD2�{!xxX�\?�]g��ƙГ�� �D�J���(�/���p+hx�x2gV�ܺ�#���-d����듆<�h�h�F7�5�6�8��QH^nr���F�=to=��p1LBaY�%\���5��,���ZY���Z윦��`s�o�h�'KA���ZwCjv�=ԵX2�� 2����7|�n^�(2�c�T��a�D������Y�S~���
]y�pӫj������s�nϭ��GXG�"*���g��v�xDk���hᦜ���W'��A�?Q�[�e!!q< ��B��mJ��ەTd��+�E����4�� ?��ʁo�0yR��C�]���T��Ի�/��1D�)������Hbe1�9���K=�\}���dj�982�ac�.�өڼ�&$ T���+���[���e���9�4�O�6{���i$�a�|��z��댄���>�:2��	r��,г�����UFn/�O�cR����8D�.�-��^U���%=�����;?��͌�
.��������=:�))d�e myԥ����j�	==���&�w.�Qd<�
D9"��"��e��WNg�d	��=�F�d�6:���u$�)}l��s!�!�le��������ʺg]Q?���A�
����ĝ���?�sb}J*��F�O٤BmQ�`�ޕ7�p��̯��w(E��9Eb�����`���E] %�㋫�F(zAŔ�A�E�;��U�n��0�!z&6�h5�'��8~�ǆU&����(�;��)C�C-��m%�wo�t��P��^R��_j��^�=s�uMaK&K'��Dj-D\H(u�j+��_�M�M<�`ȇ�D�͊ss+ҥI���Z�IhiK��]�zA���5�"�3���4�i?�6�:^-��\\;Q^}�ဳ".hu ���>8F�J\��}��(.�^�־r(=B)o���n�2wF���0<UO�my�G����!*� �i��&~���Ci��d���gf�60_�"���ҽ�A���%���H�ZX���VWW��4���i�+HҨ��a�v}roiU��͇âx�Ϗ��;�7���2";z�	^C(	�s9*ф��/����x�wa��L�3ǁ>K�����?Q��kgU䉗j���^�p:X_��/ �f����@A�;�YR^���#�I�K���.nȨ2�N
F������ȟߨ��3��k�Z��-�LI��u�\d�z�Ҡ�P ��%3F!�S��h�Μ+(�X����x����ijJ>ር��e'-����y����V�g"�X@���L���&E�'�/ذUϫ���g64�����@u�p.:�e;���s�c�IuO|2�F�_<�!I���4#19�mQ7�f�޼�?�VGV6��qV����ij���k��G�$SA���t��f��E�|�]T+.�O4�H�c�m�D%|+����T�$�,�d~~��V-�vkZ��8�z}��W�:�1Õ���л�\��#��)�3,�mO{4n��t�������o������ٶ���߁�����u~��X�$�Ѵ�l���$�u��+s9o�$���aM:����g�g��� IB���"�t�-=�j~a�edί�S��z�x�aiTZo�s�B�I�7���t^&mZ>�[Z���68W(b���๖}�/����	�Of��^��O]�x�m���������
�a�$��7�ǆPh�b��wu;��&/K�%Lʳ��M��a��5�9��gy�)T�m?���|Xf2	o�\N|T��¯t���V���t��?��vߔPL����l�`�jzE�����	YGC���9e)'�ߖ�|K89�'�`L:��l�-�'�	�&/���K¾d�%�j�kK$};��jȊu��i�ՠ���=.30���?��#�0S�SV�#�=xG?�Gw`Y�6^��T�e��Z+��fS��|`�m�`��QB\V���lP��bՄ;�i�݃�2��
@��A��`$���2ˉ�8nMß�y�3`Ax�}�_lLKA�|�r$��T]��wg�(�֔`�m�va_��G�X��u�jI��	iO�햂S�J*v�}l��T�xm�/�K~<�8}��9�T��]��d�}����_˱���A�u���y����x(�y��HQ��]��^���dɏi y1����̐W��YR��~���*�|����I\��#��>�p�K��;�-���;ۃ��|��;��������KF����L��e%E��JQo���H�9nW���ɓNi�rڧ'��
R��C�p:�7�9�zmTo^#+S��6��~
^3�����aܷ�-T�)�#������-��ykv}!���Z�bۇH�r����3��(^�����sVKq�Ai5�\MJ+��ϽM.8ݶ��VN�W3�@+��"���u�޳� W�����bD#+mc#�:�X]Q�$%��#Rpz\Em�7f:�Q~���� Y�����ߍ,�0^���]���h����I*�*��82���{h��w��G>���ϣg���^ӝ��B�j\C�V��1�4����BUMo��K���cA���'l
ۅ?d�L5"��[�ɉ��tM]g�?y��ČS�FO`q��{�T���q����9y���-�q�͠���!1�]f��Fʯ��׹(M%���a]�DuJ�^ᱢ��)��z_��Ը�J�9�wwa�t_�ڦ���6�Y�)1��b����ȍ�S�k�7)i�i Kse�1��79B_@�D�wLR�}��H��vٙ��;.��)ӆ���kck�-��eK/���iD��֌>,�0�;ۛ��m��$|]�6"JQ� ms"����PP�[��̅���Z	Җ��uC�T��K��qD�6�������B��u�^�Is��~�S^�9�J�YNFU?.�L1���R�T��V���Q��ZTK��8��>���F�n`�wD�(���)Bne{52�n����3���bF�g�T�H:���3M�����+%���J�jH=w���)��R���H��Brn�f�,��JQjI
&RT����7�Σ��Z�2%%Ti�����Ё��h��x��� 3ep����!N����3u�j�:�D7p`d�ȱ����m�QEIǹT���O�����a��~W4�ȱ��9�|��F_��Bg߬۹�~ɕH5��,+�:�4���MZ�ʛ��)y��Hg[%D�ݮUHA��O� ���^W�;�u`r?���f�C�gAk!p}K|X���d}]��UP���J�B�b����7��,���D�i�sdz��>��64U���~�'j�1o:� 
�k�om��\̰�$��<_��M���D8�=�_�.Ve��
:�7F2�Ή�YɀB���Q��+'��]#���S|�~���Y��D���nib_�(��,��� T��I���������;$�r���j.V��t�P��}�+~�K�	r��Ŕ��B��98]^[�]�U$6�MN}��M,"�=���dt~t��֍�%R8�Ve���z�t	�ܕ�d��8�`�Y�Oǖ�":Mw��8x�l^�<z
q�E����O���iiF@�Xx ��a�s��'�&�c*ޑ�n����/lhI_�'��u�.�.�鏀<�Z�k���NdB �-��;�w�6�j5��B8��ol��jcźE �Ӯri/ݺ랜
tn��MJ;��Y\�u�D�+�|�@+�9��5�}iV�;���VVf�/[qb�!rlx�=���`2�N	IuL�Q2����ă�;F ��s��x��p�]:c�gv�.���͈�e���I|l�(����P���(Bk��,EU]��yXq�EzN�ѝϕh��!P*�\ԗ�ݹ��vct��

�h!99]��~���m6�½�4ڼG������=��yӮaʵ+`p�; p�n��:�y�#�e��Q!�CQ���	[ _�g�������̍���@��e�(����wD�r�Z2��V2�?��n!f�Ϧ�\��{���O71(���'��7�g
o�£�L�j�{d���23lU�3�v��ڔ8K�� ��J��a�q>��bR�p(�5��pͻǤI^�/�d�������o��
&%�O�D^�CA�׈�a�����@]�l���F<)K==�x���0Mq��!�3��>�a�^�x9:�����m�h{0dz4ߔ��1��$��o��t=��F�I��hv�m}���3O�����ŷ�TL��a@�Wl��f�>�Q��Q�?��iƺds ��T����%-�wu%��s7��i����|�Mo^�@Lj�[[��o��@�?~�p2D�R����B���rBeC��>a!/~}r�g����Z��%���8ߞ> K�Rba��5�x�^��H�Z�e]T�ֳo�����9�{4c��䤤���|gf�����Is�9#�-,c��@WǓ��	O�>�v���,&��K�|�u����G�f�
5�I�{(%�;�fx��9W�̓Fn�$��5M��(n�%͹���qt�z����$�f���k?���%��F�=�����c˄ޱ �&U()Q���6?/W�׶Q&&�����l�xr=��D�B.����Nj3��␔�m�RD�0T3����Eg�V���j�aa��
�p^�����ө^ڪ�K1M�Bb��_��n��8�K}!���(Y�oG�g�u��I��VcH��+:6f�a��5Э��!1\����߿9��?V��S��e���f^�>6��Aʈ�M�ۘ��y�^����5~�a	us��C�WGE�_�-�*�
��J�t3t��""H����)����� �84��w����?�w�{�9�~�~���.cu=������%q�ߡ�B
�{.�7K-���x�����G�X���f�%����g�s�7Lë�`�F��I�]l�[l�2dV�f��		>�%a!PR�������K������{U��+?�S�s�iRLx�e�d��O�:vkJT���e\I�X�7U�Єmp�υؿ�!�:=?o��K��X���>��Y��*FԧXb�ā���c\��>@�v�؁���x ����kfz&���j�;��ݸ� g�^;~'��쩬,����U��?��� �zq��25l�Zn�u.Rwb������ �=WmCfn3��~�C,]�)j���x��ύ!˺��5F�ؑ��o�W�(�u�S-�O���nI|,��f�~�G��!6��t_^��E�E���r�y ��c�K��̙����qۀ��TK���O�h:W��V��#��>�b�z�׭�S#J7�_ �L����~˹t����g~3*"}]Q�]u������X �{��C�a�
���K|��3�4Gg�:� �b�]ٓ�҉���J�
1I^ܿy7&W|7q�@�R_SE���L\f5�`�;��w�\���D���̌Kar�VŻ� j�?�m��N�W��ҫ5��/��s�9q�̿�+�� կ�5��}��������`��Y}�����u4��#����l145�F�/9��o$�`�7��1�e�}ʯ��5��F������MWH7�i�~��-e}��S_I���!v����Z�@C���XUu�@C��޳�)���K�g_���7�'���W1�U���h�D]A>?kqw��`���+����e�����e�k�<�|A��r�/5����#8�I3u��/O�L���%��CAXSu��<%��x����!p�w.�3ߎ*{���nwٰ��/7��SE�������*{G���>_��
�b�sU�Yު�IP�B���R�ohW@���)P��]��WFH��"�{l�3����]��sk)Қ���ff��G�L�f�9*����[>0���80.]�7��0b~��9��U�mb�k~-��B�[_Ϫ��j����0Ng[aD�r������1�"^W9�
��_�����j9gpZ�W�K@8n(�Q�n��,�w�0�����n��G�Xz�B �T���*��֨�ycv�l�_�
V!�H��0,�O�6CJ��5Lz��e�7	
yai5��f��g(��x:P�uhp�aEC�������ϸ8;S�Wh�Hfቚ�������_8�?k�m� �Z8S����T�����ߍH7A�l�l����jN�Đ�.��RбG_�g��#�5rE?�\��k�⑸�6�i�Db�Yܤ�В.ZE^�8=���\Lw������d1�y�!�7�)�29t̂�h�!��.r�E��Whawv��K��*�8e�V�x&q��Y�`c'bl��I���Gq���s^��}���@�5�>��0�`]OQ!����`�/=�Q�r�y��/8�l~��3Iݴ8!�F�%��)d?޾��>)�[�j{�sl�_є#b�]���'wc�wR���YZ����9ۮ�#~��E�܊8;����J�M�o�h<�������;{e�q��uA1k�3��q)�����������y�`�e��'� ��ʼηͮC��]Z�ޮy3�+F�)X[?ȏ!�
9lMEmg�(�y��7| 9I���-�L�/+��y�r���@�e�I����o�^��tY��NN�}��lh���vJ�2fySb���]J9��^��x'�Bg�g�~����8��]>4����R/;:�Q�HX^�]��9eH��� 
�H��/�}����5�9�i�����	x�j
S����i�]e,��&G��4K\�RB�����fX���Sǯ��Ҙ�y��W}u�S�~���|D�a��{���F�������M�M�q{���c�zgн.���s�7"������mx/�S��&�'r�9�MM�3q�u;�������e�3�.ާ	��D(�j��[�\WA�jۥ*�ӓ+"#`��sR�7��a��������D���au���#/|���[fU7�s\<�#�I��ړ���	sd5��4���oBڤ��9��}���� �k�1$��	ǧ�Y"�k�˼|7�lAA!����2Т�S�^m���֪wu�J����&^������Q9j�ҷY�>�}�&��e���M��
�
�-ѱpIs��7/t��0V�$��޵���|�W��G��S�9��R�zh��OcċZ�J���l��D�2��'��6ɺ{�!��h�����?m�ͫ	��ddd�mE���?W��}!Qi���r/'�1���Z����;�S��?�3"⥎n;�_j�^�	A��)�:?{|����X�M��lB-����<��fU���ǽn�����������D�\��;�f\�"�o�錿�K��	T s�@����PSaUU��)�r:�A��KXt��TtY/�`\��g�M�_�|ݨ��6Z�{�������$���&��V�K�$d���r�h���Ʈ� bK�6x���~�+�+�.i|n�� ���g6G���zW>ⱂ�T��ʂ���m]��>?p4u� hl�S�ּn�k/}����?��w��{�z�-��V����Z> {��}K����i����ZKIঙ���o}����0WV��3D�mM���<�����bfa)gYX�������+M�au��Zi�.�Ĵ���/�r�v�
��0 ����E��,������h���|
��\Ϭ^/��ߎ-��2b\�e|�x��cg�fX]]�t�^��ϗ�%j�޵D���1�]G�n�G�9�RR_�X`�%X5/x�����A(��[�Z�.	�	..߾����;e��zcW�@dV�8j	�7n�"�9���FH��46��ּX~:;�,y��_G��mF�ͼ��3�{!��>�3%����]�C ��_��?�+�<��TC�ր�q��%bc�a�g���i�A7�A/���O�>���I@D'�E��ȧ��j?�I���ǆ����'ە�P�	3Izu���x,��Ŋcu��Y]���=����*Ʀ�|��P�����:	V(B��so���ޫ���@r&Ǩ E_�QN��޺x��ѝ�_Uu>�#��܈k�����,8���pfB��J�db�Z6��G�w�x;�&>,f�f�UA�IϺG�j^�wi�^[6�\h+�u=��n���`ӆ�Nϙ�q�w Zbs�>���l�Wd�K��	��{F�%vj�u0�̂��K�mQ?B �a�{�sT��x�j<"@8ʆTk(�t3��Z���U��4�������C�//��)���~�#�Z�~�,;�R�W�AQ�U�&����G�"뽸;~|������s3���5;��#L���FB�t�t{�~���2�b��ޫ��G,��ҀF�O��5V�������zn[�{I4e&�����'�5��9���EZ��Bt��@���g�7_� ���"��vĔ��CbgW��u%���*6L'M�d�<2Iu%�*W��O�=y�L�1���@��ذѥ6��qx��QX)�?m�KP�,�4�Q���|R��W�u{��{x�T�w(��Fn@��U2��ὥX���{�b--j˴�ϨD�JKg"�g����u�Y�$�_��۝/w{�eA�X�����_�����������Rw��nQ��Fّ������4y��j8�\�q	]u8����Q�#�n�����tN =½�I���˹�e"�vDY�B��(W����Y@����ZDC��]�q*��K��IgF�u/��
�6��8�P�˥��C2�Q	�=��L�'u�"͉��=B���B��f
�i*�̧�#T`�/7�k�'w%�I��&{��3���c���G���?��7�X�p�Y��<��[?�+13	a���h��\#Gs�«ĖBƁb��\Vj����D���p����K�C�1�so�G�&��FQG�D�^���:>�A�Z~��8N;+����JD��!�j=�e_}�S�����<#�#�Ǉ�c�J^R���K���+�^s�`����//1~)�����Yr���U�h��)��~Y�Y�BYD����5w�x�1����"��j.~Fw+�Ԥ�� 
;f�
��.���8����ͦ�?�L��z���3L�e�=��Γ��}1�|�{����Xj�����l;kDʁ�& )� 6���lӉ(�#�J3m]����I�o�-��0V�sWB'����CZ�v���� 4T�+�34p�Yyt��wY=X���v������8��+�u� �?W��a�闙ߞ�r����@0څ��������T-��?�x��d��S�s�ib6��+��[�y~������G���'����XU�m1�ؐ� �=�n���$/���'!�%�4�g��vȜ����va��chr\K�ZU�x�D*k��5.U���2[�?�� ��c6��Aզ$���\5T
��s�-�E�'�Q`�j��/K�� �0ܦNV2��]��ͣKe�^;E�[��^󋡯=Ml�ï�-�����Ǌ��kQ��� �Ro���L�?���u�%y�{�1]���w�?��EI춿F�ə�UuZȀ�&�Ǌ�읂~�`���,[���P��/G�ŔO%�@5�O���W��9>z�F�o��w�њ�&���	��w�`T���\_���R�.X��q`AI�eס��ػӥb��9�͙2����~j�XX*�@k��G?w�n��������\��'�s�:���Nd[)��� ��h�E_��?Z'�i�2 �.����9�5���n�8�0��,k�fᭆ�3C9�*C�=֬v��(�=����]�T"�VI���ūY��X�`sw�ƥ����G/������=��&�ɬ!��\�O[���q�2W��Y�|�4��.�"���U$�{�|�Oc`�=�]�x*'w��f �G���s�F�����m�?����ϯ��O��E���K~[x&�ra�o���r��a��y{�����Q,�u���5�6�@���%� S�o��Җ-IN���j����q4R��/�V�u]���f+��KPjU�K,�n�EJh��U7	�;�z�Ty�{eK#z�t	�am�{Y#��8.��I� ���Ɣ��E�c/v��'���������:�a�g�oԏ��!���N�>V+�����缡2C���	���jF�b/nqE�F���Xi��A��Zk�T��*-L=]�w�P�yWoC[��	f�$^��r�HF�9u�k�
��S��������������--t�j��Lm�]�Q�T#�#���z��%��Q
ں7��W�i<��Dz�4��Hh��-~�⁠�I����.�;xdD��騂�@%K����o]���j2�-��CǶ�* �ir���oKUC�<<��̨o�,�kj�����%��e���6�K`,�p�!s��ľ.�`��6�� z�f������������P��Ʒv��JY��̳�;r�gGn�Y��᝹Ej$-�ˍ�{Pj������ᆧ�D�>�ו� ���3���/J�|5p��2��ҁ�dm|��TËU��-ٓ�)��Ex����q<�}'}we�ǳ��n<����v8��a��1�~������y��U����j7��%����h��3UGT�/�: �W|x Rk5��e3�A�ŕU��;F1���@*�npN�N��Ӎ�s��hL���ޝ|Iݽ��@2��L-��
1�T�e�z>�S(��W'6:�����NO:⣽f��%�0<�g�U���;��53��V���&��W��Оp(��E>����y��"�(���^)�>�	�5�VP�3Ѿ�5$iG̞�p+����Z����$�"���*x�������n����{K��O�`�V��U�������~�n����bD��]��Ya��Ս��`��e���kpkY5P��|h���jeik�(0,z�����ݵ�6~>��M�i����?��k/>֠��m�G�[���@����/b��_�U�Ѫ����fr����ru\�Y�����w�ǋ�H��v���V��)Q���(��}йKq5���Yw�W��\�|475�b�!vtЪ��r�����R��p�OD����?�q�P��!V�;�g�v�h`��ۯw0".$=w�I$yR`�g�Jk��j���xmX�Z����47 ����l����]@z���d?��@Ϡ�����I+{J�Ҕ��Of��7�χ�rovshT_t�l|���-xN�h��'77ft��Y��y��B���ܬ���X���p����~�[�J�U����g��Ԃ {�g}�zvg.�9�t��<��c�xr>�6L��p,��D4���Gg��P@���%a�⸸��Y5���8� ���)��V��(��m�|t���KP�;��f�r`�	l�U� ����5vt4�+$��s7t�s���[��au��VȲ K��F(��H2�ֿ/A�x�gU�*q�-Q��N�~�%����N�d&`��]LybsO�')|4���Ҍ��E�����YG�ܵ�rd��DA�5?��Z!n���)I� ����s&R2(�w�"�
�`���p�PD�y_:Ŋ?�&YF��s���jk���5k����V�s�ֱ��ϟO��d��L:�''3grc�g��{KH'��»C���8�щ���͛���j�ےT�ƛB���^?�Q�2j��U�&v1C�xg]�i�7���:&�ޝJ��mq��0�0\��$������� $w��A�~�r�D��jb|�n�5] :�\3j)��X�w��xs�U�c[�7������C����ᄰ;!�!��p]*�R�����(�T �T^ԌpH�b���p�f�С����g>Z��{H�]��[�zQ�꿋_y<���G�8*�j��a�B��fi�$2����W��^�����$+-k�*]�I�2��x��c4�̂�Fϴm�}��!�c�7D����T�KN�
���&8@gn�T�%��b��i�H�er���鹍���&~�З��ݮ*SL�@{dy��!��ҡjωu�nЊ�Û?2���o�5�wtb�Y�������q�/��f�
7$���x8l�`|q�ڸ�,ps�_�dB:o �3�ǈ]AyvlNe�m;&ޙ؁S�?���͊�T����e�j^*��l�n���l��W�E!C���u��_�c���G��3��㖋sh��n,%C�~��LBI�F��b�2�&��K�����纵�n��8�*�Q�~;�:+V�c8C��3pa���!��)���â��"<1�;/�w�X�a��F.D���!��ӸD*<v������:
�J���厴1()V�HA���u�r��.���yx��-@�m�^T����t��R���ki[�]��pJ�z�ZN�����}W�Y0�ϜѼz�� Mo�@�#�U�r���$�����%��m?Ha++YR`š�/�� �w��YH�eelS�t1H�w��;�]�>X�C��Y?�dz8�o����������I�#ѷ
�a�Nw������� [��B�����	w���J�h�����B���O��	J�?���O>�5�����ؐ
��0�nL����_ItG���~�a5\Y�0��G�!����8�Y8W;�¯'�)����5;g
��A�{PtU��b����T�@q_����^�����T�I�P��,�|�b�ycYo�p�򪳹�����i'�U�l��T�h���"#��B�� ׯh;��t�ZI�;IVrsO�vU��_�u���/|������������s�8����:�Ñ�Z��\�?D��wڅ�t��ڻ궋*�xG{
�c�7�]�y�H_Hj�(�؏��,����3=��4n�����C��S��ȸtJk}1�u强s���Z9��	ph�2"6���o��Y%Jm�,)kD+wқ�:��Eh�ne�V�)�����[[���Bsq��2���yOo��|}U̯)�����T��(�S��|d3#ק i!B/U����t#�0�V�r����xA�ط�~|(�	�QG�*k�^=[h�rnk��T��
�k4�5�y|$��l�w���
��G���G�`��{L�J��y3�0����|h��i+@��ؑ_)��ۡ�#�9U*��+7�]Ÿ�)�7��IXI���7����$�ܻ����]���?��n
+�!��������Zs�ex|a*��!ajz�s���V�a���_"�U\�����T��R�qt���JW��}h��`Y|8AOjI�&��v�F}����8*�Y��8x&Cv�n�QZ�=v�{i[�0��wف�Ij�y�zUw[�l朮<L\F��
S�ڦ�"�a�hN�о�+GR'�������/��7%��v�Vn�W��ί�ID�~�8
���%�dH߅dސ5�$�����������8X6�"�������v�����J��	'��omI'�Y����K�[ m���Õ�izso6i�L�,�������3Խ]Q�meg��\�?*k[�h��z��L>���xm2:B�+�b<��Y�6���6;���m@n�,&�[��p�"�'�Aso�J ���*����(��g�3���T�o�`���M]�t����T�l�E��(J&��lu���]8�St��Ȳ7��xk�`Hm��(qnN�:�D�F|1�]�=��������/�:��M���;�;^ymz˅J��h��3�b�;`�iY�V{ <��Vek�+|[Q�����~�������9��֟$��tz��"+R2���9@`�Xy��́���ч;7f�!;[�����O}11��ļJ�<m8�-.;�	>�*Wb� �<��:nb��b�*KB@��Y݋���Lx��D�VAd�qǧ�28�$.-�S~{��a�b&��ƪ/w���~eR�����i���6CC��¶s��4�wg#�]\z�	��NN��tn��j5���λ
�S�A�@0{V�k�c�
����ԧ���u�X�ɝ��M�3��L��lf�R4���:	���8g�G�P<6��Mz���k���8><�rXس`��/P��[�0���[װ��d�>�Ϋ�֚�=W��>e�'�Fv���u�N���
�D�`y���,��M����"x��m� gp�.>lFn�����BH_�\�� $#�u�.ǱG ��ʕ�Xc_�u@���>�GMf]�6��={��B��<�|hx�~D��"��S���7��3NBR��h�,D���#�m� �&xYMZq\%ak��D�{�. ��&\�a�PM(�`v> Ř�<ݠ}�4����3�� ����Jb����4�}�=��������5a�"�����X�>�g�9��qD�{m*�>�o�/|�Z[���M4�9���Ih�Л�z7���{�㋾�F��i L.g�֠�`F&����.��6χ��>�MO<慍X�ݬ	_�g��wC,�Q���r��@�T�q}ݻYD��a�x���ӧ,nG��^^ۺ��%��o,��p��b���O���L9yk��� MRs5�i�Q<gbg�o�����(�^��}�à��'+�`=�8d�z���:鈧�<ַ��5AWO`*���o��c������r�a$�$Û������S�}0�
����%=g��LS�#K֒��?Jg�%��\gP���n��뜚��Jg5M\��Vh)�����r17p��o�]�����s��������8=�6����4�XM�m�[HB��̑ �x<F��T&����2�C�bii �TF!��;K�W��I�d�w�"�&Y��\(����exg�fyD{�p{i��]_(����4P`|�z~r+��-mB��3��~PA�y&�j�?-NUt��'g�e6��m?83%'	WS���7y�$.زˈ����SD<v/�\�QD�>�5�	2ץ�/^N�u2.��]����=%��<�砫+�ֽ7�*8�q�1�ݓ� ��Pš��d�3׃��Ҵ�k+�oަ���X8�̚�[��ȑ�4!BDc2bi�6U�e��F�0���$n��!�(��[�T&M�<s��m�����w�WM3=ݤй6��xA�)9fO a���7�OS���Wi�0f�Y���孩6uW��nYQ�`��tpgu
�����_�W^-aJv*RC����+��KL'���z���������Y�6�fw�<��Ld����@�}��=Tm�N'�VK��r-0�%��I���RJ ���g��!�z
"���C�V����H���q�����m�ū�!uv�Q�lnHV�!@�[t���s�IH;~W�&	Kij!��Va>LHUCh>OG�z+A�j⡕Fc��v�dj/F��G��)�4�$Y���L��?"�{w�۟8&@��ː��2Tw�2�h�y�����	vĈ�_籺�s�P(c��|5z�_����Y��_�6�}1�}�Z��-�]�΁���y�5�9�g��E|��{A��%�Eǒb��/��dՖ�1���0�`�[+�R)WOk=��Ց��%��C�3I���,��-qT�$->��[��eShϙ�1!�ф�օ�su�=��æ�> N 0���|j9�Ί��`�����,�s��=(0s\�%�h�=��������v+�9�Ry��%�r�����"���S�zz!�fRwb~̃�ɛ�{KD�ɶ�z����J��$S���_��D�?Xu��pr ú�s��8� BŒѶ5>:cg���ý�4Cc�.P�C���E�MnQs{�������̩4��J�Z��v��[W2�nq�[�EZu��CuȨ;y��`Yns��,���O�7Q*���V���(��j�'ts.J�@+���L˹+9%�V�nJ���Z�ۭd�S����aH��[��}��D���Cx�,��@d�wIk�O�7�^q�$��{[�反kDF �n��Z��&�R�-�!(���8�`_�|�ɛ�y!QSf�3m�{�����������K�H�(���y�����i&(���QCPeH�c��qX'��퇌���r�r}�\���
Y�ǥ�{�@`��F��qt��ַO�_���Z��
*��N�pU�C��2+�%��<�����zҮ�40��M�}�����5z���HQ�vv]%2�ށt��,��h�a�͑�+�G�:� O���J֕�K��������)�F2Gg�n5��)2���hkU�� �hfSn�����D�ߑm�@�(Eg$N�fit��v��ரn����n���~����3�5��b���h����R+s����vJ*p�M���\�J8ڟ+�8��Qwxɸ�켘#�}���1=j����[f� �$_.VG���Qm3��IK��K�{�	��Fǫ
<cS&r��9K�X>{��Y��9�9yiʁl��vvI]Ł��7�?"���p����h�5��k�6��*�:�/�ߒ����YS�eWC��꫺��؞�),���3u����I~�;�Oc����q�.oi~�Ǹ� ���!ڄ��`�a���Tmp_/\T16���@����ieO�!�c�Y�/u��o��� f3}7"��Z�ws\�#��y��=z`����ՖƝo*t���W<�W�&�ذ��X�n�d�g?����^����Ϻ���xg����Gy���p�K�4�����(��&F���j��n �}���nvia��WnI�{c�d#�p���;�[|�k�� eԑ��y��Kv���s�����]3����\����5��]z�:��:�o�b�B
;�sbڤJ�6����u���v��BY��z#B�zXJb�qUJ�tC4�`C��m��F7��;���;[�o�{�$�S~�8�+_�� "D0�N��C�Ū�E��3O��_��i�������q鳛rW�?g�q���g����4d7��d,��rΑQtz�6��Ҽ\#��Uw��2/���t#�.���\�T`2W����m\�͂^jeP�A'�!|��gbt�ۚ�y�Mse!�l/���x4���_8�}G"�+x���Wh"C��j*i��5ټbX
!�o��WY�od3���,�Dۛ�����k5��s[3 
�tCIk�����6�5�
�[S[�ݡ��sؚ��n�a��������� ��'����d��ދ���X���K�ϋ��(|�o�	��������
���܃؅�\���3�m��{�ra��"�����9r��tF�Q��ш�rR	�����q��|C������u��Fя$����@�Y0��2d���y�|n1w�tֹ�Wߠ�L�dז��@���K�m�@׌����	�bXqG:,�S�4z*3�*�}��wa��|�p�m�����-���&����~�x��Y�7��}���d� ����_��#�����d37�ޞ_6>��qa4��<���/�ܫ%J?ku�%�Ϣ���n:C�h�S���#�1�_w��{W�,Xd������fd�H�o�ȅW��܆�0!Ȉ�ؙ��o��$��GV�΁D ޵K�|;{�N�����	�W�{��}M;UH_�LO!H㉩�0�[��F�zS�e�a ��G����#jJa�=��nc�=�EE�}!�`uՒ�ZA��<Ȏ�)�����[�����va�NV���rl*�B*9Ӷ�B�L�r��p| ��JE-��~�mN�ѓ.�\���|�[�|�-���T��.
S��M>������ZΓ�_c-2���|Ad��w_��3��u��W���q�j仠�����42߮�<�S���;�.A���5�I���~d��ɼ�`���1e��-�K�����P����pNՁ �������!.���6#����⋈�����I��i��nI�--lېpI]����t=;C�������[_ע���s���!��4�ic��,�d@�P���pؼ�W'h�o�֝���dp3�v	�邀&�����?��% �z�4�ƃg�3�v؄죨��%�E���%ZB��2�3�G���&4|ѷ��B���9��ۋ�]IE�M�e����>�-7� �YM���\���$|�#G�k��D�o��;�o�Ȣ!��Ѳ懲��#�Z���.Qz���{�F�&k��}������wA��۵��V�m��P���X����B���?9�)U�E�E]?��xuB�5P"2F+5n�+(j�Q����]^�̅-�s�Zcixҿ]����^�e��qi͇�x�R���Ը�Nc�gz���,+�v�9N��_��-~���Dd�g�s͛\����G�۷�}J�6����#��e.�Jo�}�ɍ���7tgty)�k�)Q��_H�T�P���������N�-׼�.ק"�n�0}7�6<��T���������te���ǵ�#W�y�n跛B�
~5q@(�-o�t���@���-��Q=O�u�N�yMn|������u�1)N씅M�ᓼP��\��^�q�'�����C�2މ�������A<��f��$E�A���!�f�[�9�A��Ø���_@�������_�z�7�z��k�km�nHy�{wH]˜���P%~��[�Ɵ�	f�җMŵv$�.F���B^� 
�>l�j~�1�8�(NL��㌼뤥��=�YA���td��Jes������<�G?k��8��B���x�}�إsGcY�[?J~����G�
��ߟA83��X6w���C�+u�nc\���H�]��[�Z��Y#/n�+.$�T�{�0n�;��
���f��r��|o����kU�/��m]�9o�}�E-�^�'���8�َ�1♯8Y��߂���U��G����S -�nS���*@�����;P_�^77��2�9�^�e����I(���$u�S;�j���b�m��r�(u#�,a�"q>�!�ja?۞{w=�W��AT�njPm� hH�j��̿�(F������/����G'��|Ji�IN��MiLƴ챷�a�PY��>��'	H��/�<,�{�v�sm0��%�&����U*]�>v��-����\5[5%�w����&�����KX�/~�@�$����G/ɿ��2n?:[����4á�O���K�q=�g�l���(���CS���O�72L��]ң��Lj�"1�_7^`���B'~6[��vֱ�.9ނR�f^>�4-��1=����u��䀿�a��.��Bē�8 N��گ�����+���f��v�{�i��}�Y"��i�1�v�[�@O��S�2	��к$rX����\n:l�@�%tTy$Qmv�b�g1��s��L�����˧ܻ��R���>�׈KZ.��y�3��yMl[���Em@F��qQ�8h'}xB.ޞ�X/;z� �ڄn���r�	���]o��$�����Ց��~�@X�=)N�� ?0�	"I�����E��M�ˉj�1ŘT��+m7l>��|>�"���-`*�����m�i���h��T�FWgj�̊64-^z5'�Z������1�*5t������zb�?����^�o'�r[�vꮹ�~�w�ƒ'��mp#�U�%L|*M������I�?�1�%��?Tyz�̣�R{��cN@�w�Dq��+��%ɚ�8�K2���b��s:q�B#�-Բ�_�t�weU>��"�����?rO>��}-o�q��?�ΜA�:�2�WwƻO����Y��Iw=��IV~�\��.<d*}B1$�ٸ��#vr'<a���g���w/��+�Y�{���/�Y	�4,xڇ6Mը��<���R��X}b"�~��4U���a��N����2A ��E�� a���*�� �D����Յ8B;��*X�i�FO����íy��ݙ��H6N/�%�B��}�z��r�0�r`ɤ�������L����q�ߠG��-5ɝB~yD?�(�k3]�g�DnEx=���Ǭ/��2~���E�ffm������+ؐp�����P� 0��;�Q?�[1�z~�޳�q,��տ�{k9��Ʒ���*Ӣ�k�������E��5�ӱ��0�����s��+b��:���N�h��K�Q�^��Jq��~̇�N��Gĭi�!.�e�w��2g��ܽ�m�~xTp>�S�&uG�;�l:��x�~fTB�]Ci_3Ͽ�{���]�2s�괘��D�5���x��>ޗw�cU�]�!�R�Ԥ�?Ok-İM&���{��=�!��NF��H�����m �@���J��C�Y�s�̏�<`Dw�Ct��aJ�%�yP��
���"9�]����Ԙ����Cݕ3��}�f��� ����Đ��Ͽ���J�Z��;E�^�҅�$9_��m9�y�G��Sa]���́4m���&��c�V]��<n��s�uXլ�?W�b�X�aҎ�|H� ����8�d�Abg�FƸļ)���(�F{H����#/�=.�����
�˦� z8Wv� �V'�� GYF���i9�W"?�����C:�w�p/�U�"�D}�.�qZ��A5�A�v����K��AF �V���iP����P�UA���j�	8Š��.b��r������M�a��q�Nk5"��>/����2��㷀\^S��������CӾ|�r�ӧl����^�l~���'��H����#8nSV���#�	����4�Ao�b?�����\ǣ�i��O0D(��<���ɉ.&\������B��.�/�	��&�O=��z�u�s�V����i�U�Js�����O�������В�O�� ��q=E߯��j���������)���M@����7Ïc��,^Q�	�fta��5?_��ප@e6,��,��X�P��_t-^c��T��^�E���(|0�K#��,x�������ǃ2�4)��\oz�j�]�d���ŕކ�n���p�qK�պ�������=���/�5�ɛ{>����(ǳ<}?h��h����w⽻��㴜�\��^B�2�ã��c�/��l���X��G	Ɋ1Gn����F��kM}y��]E�!�����6��`�}��I"��>I����(N���Xrgi��O�m���R�>�y�M��>���3n�.h�	yb���˦�=J�6�j�m���53����ZE�fv�����M�t�aA#�􅀄��Ƶ+`E�$�y\��I�S���u�T/=Qi�#���v}����r��}��顸�����҆D����y��[���'��A��t��,�ˤ[�d�f�0�����tչM���m��2�5��D��1��am�A��(�����)������R�������݂�s�9�w��#O��&������ɸ$o���fL��=�枕�	d��dDӇ�%~�˷��ͼ�CJ���b(�R�ug��ynO�_+pyZ9��0!r�C1���`=��Y����'�������z�U~����Po��!WL����=�<M�6u[�!a�q)��|�6���n?�9�]�x,����r��2|_����}��7��4|G�^�״i��o�8/f#p;��God$�� ��)���*���"�9p7��)�Iif�w>���"Z�U�����C���2�۶���3���m��e��$�;���ԗ�0����!{v�`<������ې��,1="9|$�������H�JGD?F�������÷ׇ*�Y�Aa�=	_�z!_�m�$+���-[J��ٴ�>(@��F�c�NG�AH@��
]s��,�.�)�s
�V�c�7�����jt��j���*�Y��EEx���.r�pGX6'��Lt����=�|��B�}�j�\�{���̋�����m�44�ǜ�F@��E9:��&"�ȱ���n@�%�V���e��:!�O����.��`�й�S��0q�
Ehf��u�C�F�zXU��K�1�EW��G�>��H���G~����fb���ۏ� .�6��^�;���u~��=��]��#�/��BI�O��>W�E�m�\1����G���~
c0]~��{E�~����T�.��NhF,c�J��[��J��c�	�F=�ڋ��}8�mѿ�XC��)�>R½��.�.P`�:RM����,���U6[|G�n��j�94~��V����Y�c~��p��9�f��� ���H0�u�C%	�96m=��2]_�m�Z���R4L�zbp�gOަ��V��uS2<l�Ճ�1p�|<hO��i���i����<�Ɩ�4ɇ� /��p�̞Y�Q�{��6�!A�6�9ﱊ�I��������|̛�ȋ��,�6^��I$@�)n�5��x>#a8�KF4�Ͷ��O�n�N��0�m���{�W#�Jᩤu���R"hc0�(t,K�"E���zb���֮c�n�f�ׄ��8yUTœ)�-��<��l� �Ǻ��A����	�s�"�����1~zsk��Z��f�l��yk�����<v LO���+��[�iݖ��6� ��o�L����y��߸=Z#.I�u>�Gux~�b�"��`��v�l}�J�"�vJq?��[ u���&T�-]	;̕lzWX0��A�a���*?�$ i;��)�[����^���#zM��>���W�5�'���q,��{m��T���3����E���Պg�Yx��:P'Y[��QNy �ytp��2���l�/wW .��*�ɲy�X���ɲ�"S�j���^C��g�k�{J�ާV]j!�tib�[�T�X�F��Ì#��%����>�\� �7����7a��8���A�K;����~��'��Ed�>�+�������Fa�u��.�B;��9q1ra������b���)�=��Q�я?�#i���V,�XdT��4���Md;D#y_?���a|�t !q~U.�\�lM�=%DU��3�h�G��
�s���K��,wg�R��tp��#�(Xt��<}���6����m|d����Ɲ9�S�D ��we��6�Ey���6Wf���6���D$���Z���5��6
+	��h�
ej�Wkm.�hᑉk�O䍰����;_wlI��sN�[���k1Y�	�"Q�Y��A�C~S����>���Yoe9 ��|?) ���w��]��ח��v#M��3oJ�\h�Q�c�:��c�b\ܟ��SJ�Y�Ͼ���?y:��Ct6w"��� "�����J=��mbwv����#��o|^�hj��ɼe&1�A?V�+6�'���h�\�a�����ôMWD�녷"�.5ߒ����+�4��ZY(/0���_6
p�)
���p+�h�ߜ�N��Q�䵲Y��g�w���5�=$������L���"�nu�r��5�m�nE�M����z�SW�"���	ܧ��3l��[�X�r2���ܜ��F���O�X��mG���?O����^yõ�l{q7��B��)Ѝ{�۝�/x��ư2�Z�}�� i�|۠��i���\�xUn7�񜜼���c���� g��8�)�����a�q���3���)�?�l� �r�,Z���ԝ�ř��W4���
���P���+x�uJ�*�l߷��]q!U�f�S�T�v��h�6:��i>`���s��(7��˽�z�!5l�CS*�"��轗ް��M���R��ŗ�M�,'8(��/�.��&����탃����K����.�}��m�����f`���t���I�eyY���2��Bq錙q�=e�.��*�N\���=�1�:RyXܙ�]ϙ�#��o�Gx����ڐ��w�����j��:�j`朋�{��4�N�gs�јa�W�{�CNA�E-�Ȧ���y��O��&��#�3{�ҷ�{*��.__�c�0w+�J��=Fq��)�i�D���`����`�� Y=�����Q�?�O9�v�8+SJ3ߕ�۩籑%����z�Y�{�9�K����2 5�}�pP���������7[�c�c��O�%���s51�C U0#P�`�QU��D�~���s�������!���?�D�9ʵ2�0�v�&�,x���_Z�Ӽ� �&�"���ʀ��w�M>Y�$l6���{SAm���<�On��|�Gi�,�{M.�*�x��խ��7��I[��U!�mL�D�0��S�{�"F��#R\糸q��OG�d1�rj6�Qj ?BS���!�f�7*I@i�^_����KVG��8��Ј�O�\aX�v�b�W)R�.'�N�4�ް�g���$:�d>6U�y1�=lq����c�Û]�{F�	����X�L�u8 �&0�=�VN\��ǖ�-c�K{��r?��E�ᖼz]��-T���ڽ�њ��I$�����d�#��~U	��������`o�! \�E�-+=�_��N|v����5>�{�|��R#�c���R�M�K�D[g���YZ���J��w��|�v_���?�^���9���o���"�:�&���9F�h���q���Of+o�M���YѤ�'ev�W�k�[�2٠?����G��HU21��GG����[p1^���(ٱ��LI�=!�S�t��*��ru��9G�dZu��],����}��5@"�k�f3y���[>�]���P�wk�X����4d� �\i0ҭ\�u��J�	�u��H>8ݡJX$���x����,A)*O��:�*���%�)l����6�/���棇,
?�q}8UɠT���@��;�>g�1�m%��V�.]�.ڄ��@C���͗��l^K��[iī�3��V�=�.q8�US���<� �u�hb�a-:��z��.��v��� t�#�=�k09sc�{!�S�ދԱm{�l���T��p%X�*ޡ��I�I���+�y�r��B{�~A�woV�H�;OΣ�`�
p�B���⨺3O��pg!kɳ�KEо'�L�>eIG7�� �3����N�3X�����������)]Dzic���`�԰a��؞W�ı��5H������,���p��LK�_�Ƹ��4��)C�st
SW�?���zr�����V�q��&1�?~��袓��m~���#�q��(�0����uM��A�n z��+���Q�6���J@��G@"�!�
g����;���o
u<�L�� ���}��{��
�`w^B-m�ikB��b�Xr��R?�h	���j���W5#InOG&&_1W�xSG�r��_���=GNն�@=��e�~=QŇ��F�=�D�� vH^Bd:���<=��(2=ȭT5.����-��!��L�u밚�"h�ݬ����_�7��@��x��k�
,p;�E�p�xt^].>* ��h��O�]��=؃�'3q��� �Ь�{�rBH�i�6�
t��Vsӡ��~q��L�8&���"�#՜�E-�����������p��A����-�HF���e��/�#Œ�R㷲r���p<x�������������%�?�(�1�B&}r^�l�G�Kuw�z�I��OxPt7�N�$Q�*2"�z2_"������Jz?͇}�@�;Gbډ�T�8r�/ڰ;99}��v^��󼝋�h����2������Ϧ�knn����Wr{`�n��OLq*#At��(��-/�<�,ը ��$�����^�Ί�6i�������.��mW���S��+����<}��-��1�����e,v����'��]��Rr����k�m���ז����I=���=A=��I!P�[Dr�#!�>��:�<���P����K�}l�<
!ȵ��uH��9���tյn�����{L���?Y\�� F�
w��Y���B�('�ES�K>9K��p���~A{"Gd�?��7K� U��_6�)R�!Q� ˼ Q6����{�!����:��!k�S��0��l���j$��h��Aɓ�bD�swwoQP���BA���>�8�uz��ZuW�p������o��hs-����KK����/��ʍd�<c��]������)���p��h���0��:����q95�sR��NQ��E�l���ܑ>�_������
::�����J��ڥ�k�����(,"�|jr�O��TM+��\�J�i�2)$޲B�3fXL��v6�����lM"�O��3���g&�a�s�t:�:ҷ]$Գ{ e��r��E��n����gw�}NG���ew���Uݪ� �K��Kr���e���D!է;_���ȥ�#a�؀@�b��~�r�?��1(A�}���67���,8���U%��N�H���׳7V����XM�`��`��� ��A�'̜�)R˥d����۽x��Ѽ�u7^:t�r���2��
��W�%�s��*���ǋ�F.v'�IÉ/�.e���mkW�F5�c���p<~&�!O;��5Y10y������
��8RP���E)�Np��,J�딲v����Y��(�c��1N��m��_;/'���ƉY�M�R�s��dQ�Y�zr,ޠyIw7�v��o�Ӎ?��(��lup�*��Rb$X0^/�:N5��H���
�ʑ�j��/�:6�� v���A�`/v#T�',���^�3|��YB_'�GԵ�(8�?��m�O��)�+�0��[��J-~tW2mH�o�4��Tk��|�ݏ�+#��z��G�F�uC�Xz���]#���OMjmM�����w*��b�4Ǎc��T����Ō)0ݛ|~w�6��mP�,��JOo��	��sP�6���<���}Q�(v�F�CT�W���V�o�m$W��Y�
{�?\�S��F�����SI��r����j��䚽!��?��~2�^��A��1%�����z����a��?��z'f(!&m�2�k̫�'o��YM�X*b��uu�K��Q]��M�JVyypI8�Lܺ6��ʏwp7��L[��na~����(�vx<����Yx�v߲����jZc�z;��R]��L�h"����/s�gfa�����u�ؾy\�kӨ.n�E\n�m�ut�M��H)�h� Q���A�a����d����@�IY�<6��i��]� g���4h<~�Y��vvSp^R���r�S��_���_��l�E1��Y�-��R��_���r��ՃOx~�c��y�v����:�|�?s�s{Z�.7(�PfX�Q�;�d{�����ıK����iw'-wq�?�Ѓ�x���N�p����3-\�%a�x<J	�Ջň��
�d��:�|{P��2~���dW�߸����}�*iD^K:oO�D'h__����I�G�����_ߺ�2���@�p�;�ښ���S�O�W�ު\A f���F C�~�.��vH)�zS�x����7�_�0�pى� O,�u�*.���}������s�����ت~���j&c׆��x*�|�Q�>z),���ϕE�E��1�**!��zgݗ
 ��7u�Y����g�f��wI�@aK�Sƻ�� ��4"�"8^ޡ�����Uܴ��)�"�*� �]��o<4az������B����,�FoTCDY\���+�b[��'(��	�i��h6�g��pP��~c�}�Q�h2 ���)���~!ʇ�a�t9��~����L PZ\ϙ�TTp�4��X�G�~�^q}��Q��Lޞ���$804��+=�*�Q�	�q�5vJt���{�
UxK�H<N�P���Ǌ���7���PZ�fYդ�����w;6��Q��ޣM�-o��K�=�[�fv�X�u���,ݚ�ptE���wD%~ �����"=3��	#���X��GBs���S��B�ӉS��AE�>v�4�\��-5�dU\�Q�iW8q�㟁��X�
��_�݅A�l4�����y��뗢)������Z�ғEdjF�[�<�/o��A����0ȇ
�w�!k�תߠYQ�R�������P9&���<7NQ
�eiɥ��X�Tc��Íz3�_�Eb�ר!י�7��s����X|(R#����r�w��x0��� ,��܀�g9�f���5�0��C����<�Z]nz1��t�c\U����R��%C3��Yf�l�i�<����Cc���I������~��=f����3b��I���?ߋ����M�j�ZA���ʞ}�(��C�w~1O��J�C�uK�?��ªY����>̆���9��!d����ۣ�H)F
ʙ
Y׋�;/A�D����()�$�(���F��C}�h�J�9ě��<��,,����h���'��������_�oZ���*
�t{�>��Zu�;0@׏��Վ���1���)&��r:���A�[����p����~A�@�Fx�\��R�(���:��=Y^���T�UP���g�ù?�
�p-B �^�3�����7��\�>{ŋSs!x�=�z���J�f���^kDjc�l-����gk��Ör��8:���k6޽]m@�O�n��E��*�4�D���X��k����?&#�����`��y=V�핰�8�lP�@�a\�oRF��v�(0���ì�����7�Ϩ@����C�m�w����[xo���`�p(��=m{?&��qf�iUw��T�Xݫ�xm�E�O�Y�'/���=�k���㿽��U��3[+�'mm�`�E�����	]�ZiW_�����Y��r��M���-s�-o݌�:�s#}��z�Z��N���� 4�霟;]n���E*4lht�Q��}f���7iwJ��n�3��D1�'�a[��di���E9u����װA���
:އ���9��lWN�`2�y��@?�_B�%�pc��b�X�e�5�F�K
,c.��{ yl8ٚ@9�ߞ�Ӧ�����t)x�z�wZmW��W�.ۿ�٫Z����^>rS`<-�a�͋���K�|�^::�A�/�HZ�W9�y�*������Ye��<�ޠw�)����!��s%��a�\��<
�m_��RK�j�+�U�՞�6Hp�-�o��x��Y@m��-����Ѹ��%��ANd���!"��(Q���Q�X^�ѯ:x:��`&���"�w���b�}��9a'�ɥ�!���D�U/�v�x%��ԓ�g844���s��~I[SZܜ����_���b1{!9$,�9L�x~�*f�Kr�A�z�t�)i44���[SWJ�%O��J�R����®�e=I���F7�*~~d�=�ֱi �]�t]*���ҵ�l������c��C��h�@�s	-Y���=��T�J����/G�~g��wcӕ�D��t�ױŻ~�~���e��K���#��Y��1��j�x��m����a�c5#����1�g�a ֥./TYjLy�|�"l��~z�w��"��4��k���Y���bs�/���{˴s$��[��0�H�d��-�p��{BW_��wK�O9�^��y�A��E��g��6�TY��o,�Jt/Ȃ��'�?��6%u۴U���3�/3܅�gm^.�R� �/"�Af`���K���/8��p�"�c�p�cL�keiщ��1�P�x�N�Ag�A�%o}��3���!����D�����J)�i�����U�I���;*v�R�)�SU��p��7>��u�w\\o"}�Bi��0� ���c��P8���v�c!c�.*h~�=%���6;??�����ʯ0��Po�o���\R��gB\_ ���< �ag&_IA��=�}t���<?�ߧ���[zU<�R1ɗC���/�������H~��d��D��Ie�M���6`*�TrB��bkWJ&�R�����:=�Y۽�х�W���^*�^����"�[ qʀ��WJv}&صuVz��r�-�Tr�v��d�>[QЁ{��L!�6�/���ܼM��M UŦK�Ʋ6vU�����o�B{{� ���Bك�������Ba��������j���ik𻦯�������Өj��ݘ�uCZ���Fg?�g
�������.�P#���' �����T�"O5+յ=F�bf�7�T��/�n�����(M��b^)�m66vhz5�����?$���1S|�O\2�3�7\��տ)�kwнUjO9V#&CTH�,�C���hw<� A�&�_�%E���XOҡ8����������="4����@]�e����b��LV�����xP�6m��'Nk�����$�'W��}A����"��6w��z�ZJw  g���j��py![i�����8����t.r�����1� �vq$L�`xx���z`�甑[��ї�;HN��Ώ&M��:�K!��ho�����w�i��/:��x~M���I4��:r�H������a�|��x��D�/NT�n3t����a���陯=���i�ߋM ���,ڸ3v��~�(��A�F�h���`;vm�.%ܕ(Ur� Y�S�#b��^�V%�H�WL�r�����fk�H�'c5)��:�/-�]?�Gz):�B�%<�<V�9�W�7ߝJ�%�miu�F7��O��N.}TĞ ���E�-%��v�����mZ���`5
#�QV1XJ���|�'H6�?����}�5��8T#�q����ό�B��E;*
��3�ئ����6�� �=@k�r:}�n1S!P�"7���H�x�-��a9T�i!u���ȳ�3ag��%re������vMcj��D��+ ��=��J���w�wo���[�.�ݩ/\蓏ّа@.���vww��M�����ȸ����oz\�Q�x,��t�Z$V\2~s�m7b:���T��¯�>8:��]�j�Ѷ'���	:�f�U�93�Po�rzr��,�� &7�"�!Ck�@f�R¿#��UL��SU�f��A��@jZ��قR��ч� �
a�@�M�5���;ྴTѮ�W�k�:��d*�wT�N�*��#\�0�]ɆJ��Y	2hk�@�Y�}+��V�8���X ~1(
��ЉR#O����+1fw��ˁ�qZG[���{N�i@7�����q���bU�qe���6,�H駭�2�\*�G)?䒦=�6��ho�4��,�1/#�v�|s�h�W�priG��!�k�"��g(�
�+6��L�L����p5�X?�#'��Bx�c7�us/ak�u�S�M.yu�v���+��Y�37�j��ħ^G�m�wm����N0,HdH,ҔOu��Km�p�����)��w#��(d$�p��^�����ȼø�9��!�KV~}�|�����bM�#�&kC�fn���~����|�����.)M�"���U�Z`ט*��Z���$� rP6��(*�GM@+]�//���(u,fk-H��P�X�cP�T&�<>���ϐ�2��1�w��
`��U�~�y�����@�<.��� ��ׯP�<|s�D�T��%!�_��#��l�#P�N�dxp�㙴�
g<~Xŕ-��-"��Fa�r�
��N�ճ5QV���DǨ�=b���h+��:��m�ɼ-��꥾��9j-�L� �F�<��c����� GC�؜���x�u¥�My��|5�W;�uwL��&�K�j����/�֚t�gˢk[=T��BB�����H����·_��m�OOO_"d����vzOz��۶�E�tsɠ�Q�W]��/�J~ȥᵨKW���e$ɑm/w7/͗D�� A��3z������H�����?Z�\�����c�l��Z~}��9�Z�P������%��"����!iٯ]����׭�K%��%�F�#��~i���������>��<�Bվdz���TO��J>��&�s���>4���y�/>
����L�?1.FT�p"Z"g����4'̡�N�-vz�g����y�Z�:H���]	�;kD�����V:'�3��@p�	} �``�9��J�#A*Vf���,�k�U�*���e�R���]����=;�B`~����"��Y
��]��qjC},�U��D�8:�l��̲z�zn���݉sʔ�I��������X|�$χ��Ş*r'E�	)���[H��ƈ�-�J���+�9�m�z�t�VM�0������:k��{��h%ߨZ�kE�ŤK�o:��k�p�R>�[����=���U&�=Â�bnH��L�-�R�8���,��ǫ��E܃o�-��^2�\B�p�D��0����+Q��ź�`6G8�m�3x_� �.n�э�BƮˎ坟>q��>`v6y�y��8x�L�n�Y3�RБ� �<|q�b+lv5��x��|�'�>̈́��S�<Q"�4�[��Hض�!
���]a��P����!X�����s?1C}R����*t8g��W;�1�8'r6��o�T'��{5���B$O�����@������$�/򾟶��n�W�$�R�V�$�ܛ�^���o��]��n_�(y��kZ
︰f �o�`FϻW}3�>��l�c�`b����Y�� }~z>$a!v��+n�g�-p���$ʌ96��0M�$Zb�J'�5�j�I&��R��1·�^?���R2�bd��.�������������m�t���%P�UH�"�~�$�����ˀ�Z�xY�j[��^�]���X�kS�v���b��ÙV랒ǘ����0#ˤ���)�PTW���� �ew��a~e&ހ��5�%�z��B1h�o�<�o!���-ګ9R񩁏�1.Izy�9�/L���}ǧb��|~F?��d�V�=�#�!�o�xޓ�C�c�����<������~�!�A�^��@�q(�0���p��Hs����擑���/*do~���^l8����H;u`<� =��� ������ȭ��W���
�v���qƢݼ���n�0T�8(`TU%�Iv�{��ǩ�,.��c_��3����UC!�#�@!���^�#��di�=T��d�7g\��ܾ�߰����c@��c���[ጌ&5�#�9���L��Gw=�U4������]�c��ŋeōY�k��f����Ee��*����Xm�6`��K���HĪ���Պ�P�p-K�{��K4ȉb�%���q ^�l���C[.��}~�#���'�^	��_�Lk�DY��wV:=E^@�S�M0���[K���U�%Ȗ����qL��OH�� =�z�R�W*u�_=#��fɇ�a��GRSs�K6�IO�7L�ΐ�����'1�Fod�˰�67���?�0�&�񪪫�]�TK"�Gx�x�XaY�\*0��˿Vʟ��b��9j�j�m!�O�����j;Q�E'����d;8���<Z�vO��KṴ�zdG;��+��)?��)0)h[BJ������>�.���j2��튀|6\�$j �@���F�N���82X��nG��W���.f�@W�l��f��[pY:��m�D�v_�*5���r䁱}�|��@�_Cw/�
���3�����@��ViZ%Ѩ[TW3���i���y�^_��⻮pCv-��{-U9� ��N�=�[�z����4`�щ(��g��%��g
�5v/��h��V��)��E�53f��On&s����gx�PI�U��sP�V����&g��l������Z�fR�#g(��¾�[��*b,/��5����r������y}���f,ڦ[F��znj�������i)ua�ٓG�G8�>�|��F����!�K"��\����9�~!�`���� 	�]Ͳr�l@�8.w���{��|��i+d�Z�Dm�!,��V�U�~.I�(7�K�������|u�i��ؾ��i�sdѤuu����s=�����Ts��1m9ͻ��e�"h���b�t3@�m6�j��}#��,H�<�$��yx5�$�����(�j�US�	VM�	���r@�Zp��	Z �*mE��4��?���Taim��]ؿ;�g�Y�� KFrux%A���I;j��6c�\�Q�R1tH+��q1ql��Grm�1�T��el�f��KO;}��i��bd��CWe}.�A��=c��́'��N	!X��sm�o^�����i8k!W�Hډ���=�x�}l�إf\;�w�S,3/\0�҂�SZ2'���-}�]�7/ٛ1C�ގJ�(Ĩ�(��)))XX�ٵ&fw��Q}���!"h,	�t��H��?� ��Og��m��9�WJ]9Y�Ҵ&�o=T��@+M參$PoU++�pv�7oUj{yh�-�J��p����O䨨������o��~*K��q�w������Y�|Ŀ*��*���j̠�hY��s<����֎�W��/���G_H�6���o��r��ġ�9�>���1��V:�5��a����Rb�H`c��"�/�T4r��$-k�œ�vy�L9�M����T���t8�Ӫ�{8���ڢ ���m�b/%�
��#jv}h�-�A!�/�Z��P����4�	�[�r1������e	��o�,Z
:��+��5 >�#��؂����=����@�O��M����Vȋ��iyO�j�Y�����u���`|'۾A�J���Ʃ�f�i��k�����������C��ï]eQ��S��i�(ť���dL��U%����s&�
x������X��a��	��x p���{�34�:&ҕJ�M�~��+�wyX�� Ny�D?֘-A�Q?|N�{q��X�{�v��W��yû�?_�?t7h�Sl�1qr�!�B'�o��G��S�^\��J5t�]G	\� �����Z��A����(ÿk=؍.Uf`p�2q� �1�������p�_��Ar}dk�_=<EܳC��S���
%��u���'���Kӛq�a#���7`@*��\*`��ޱ��9�
��p}�F�t��an^\b��{��k �e
�z'v:0O��e�zIZ�%(��ZF�j��[�b�-���qp�i��1�}��H���GbfJf�c\L�?�Sz7����T3�fI;f�������27$�m�Jp Zpe��~�������<��zY1ƞ��3��=r)���X��"�:����fƵd�e�܈�tk���6b3.���5E��2O�d1;��a�?=��j�?s��W�Zx`����)L'�c��,�?@�?�S�'�j$sШRka�<o�R`�������������z�A@=,Q"�5��FSA��z}�)�})NJ�����ӵ�鵌���HZK�ps"O���寤]h�ꜚ��e�:�Dե��7����>t������?�⬃s�Z�.ڕN7�d(K�-1.�L��!����ļ-�(�GD�/?���>������(K��b��ag�4�Q���X/�T���I�t�%�=zA��*��"��2`P	��6v�tf�/�.c�a����S�Vy;-H4q��9��` ,u����G"y��2�T��V%J�����EW����*�M�3��k�m��l��i��r�8&����u��x.涆��:�>S�`�]�����U�,i�ȝ��d\��XOyb�����t�|�Z����ʣk��3��I��+C� ��	�Da<f,���}�*�:{%,~��ؙk�mF�J��t���mry�ˮ�L�B@]T_���0�ه7Y�|O�5D}"��55��ts1�J���!"�f$�ؼ�]e��*RLC�QH���O�1��gD��,�װr��|��c���ۇg�ӥ���ʵ�Y.�צ�%�:��(�Q%;x���m�Bh�s��SN�b5�L���1E��؈p^F��W%��x>[8t���A�t��"ĉ����n����I��a��9�񩈿�_�]���(�x��Zql7e�2
D�����6�6����-y�).7&��u"����T^\��N�:��+ѓ��6����=#���JVm:�3�"��G����y�8h����6��EHM����̟��"`2�{���w"���ϼPw�)M6p�6�G��On�f���`��
I���y�V��7 �S��=;�/O
���3
�����=6f�`AY A�2�I��ˤ/�DQH�*��+b3,	��)rS2l��2ߺ)|�L��W�)N���]���j��g{%��Sd�0���B�6�~J��8�	������w턌&-�����`G�uf�E�D���:̡�A�J�`p$�.��k�K��Oo�>�{҇�f˔�e�ڲ�a��Y�^�gb�����|m�Q���1I�g��+��h盘QU�e`2gHFE�9�p�-B�x�� ��S�͋�A#}]���::��׍�H����$�u����S�q�@���r?у�g�,q��v��w6���Ցk��Đ�ܦW���ׄe�c�k/ڭ|}7�����������x��cnRL~�,�0�3�O�6�)k�!�L5ۺ_ܽת���h�VB�9e��!p��"��&Xq�o�m��xAL��r�1���P|1��^��q=�G��nS�<�;��Q5���۟ݝn���y�k{����d%��kJ1����F�]q�/��z���-�n��[����n����9�o$*Qo�����<���#m�4����]�4�c2e�N1m�(r��|���o�b�}V2��X�ͅ��(��܁-+�Y�=��ybb��]o������𖀗z�Epi+�gV�h�F�VلB�`�59Z4,�	TuL������M�9�׏�������}�r�2������;�ܥ�n�f����v�:V�TFf�r��U0�{��yb�K�g��=(���	qw_},IZ����5N���e��s[��Y�3F����&�R�~�s�����ubۭB�v.�D\�#N�����Nng�A���~C�_RŦ`�9B�yt��ueX-7nz�؊��*���͖7����u,�_��|�c�^�h2���7�Ե`��po�BD��i��s-iM�-����t���QE���G^2B%���$��ё�T˒��	���C3��So��V�VƷn,;|�T#%�i��k5����.��M�q`cC��q��#�1���&��<3D-T1 ��8zp�'A��Pʠ���;f�&0��ƛ�+6>	�Bl�[-{Q�J�򧂷�P3���¦7;`��o�Sk��0�(���$&X����Pݼr��w^��(ή8Sy�K���X��O�z71Y��@��5�Q{�Y���Z�ҝ�B��҂���d�����9��=�ve�5F�o~*���9�3���sv�<7�YBl�~�=��pT��cz��CS���$vp��T�n��8���H��7ק$�\�����8�h�Ed��>I*l�K�s���9�#������(�����g'��Ĝ��{��{�xr*^��/N���(��'��K�q9�m�9���.{�3�nN>��cGD]�s�O}j��:҃=Æa�Od����f㼠��Vw�MG�C��t��1���O�����Q���ϼ�Sc�?����B�T6>l�gۑ���Kf�<��Tv�@�vo��gQ�����"f������sͦM��(=
R�ȵ��/�]�V��˯�$��a��K�Y6D��a,�,�i��pby�m���(�1�����B���%W�KJ�2?���wX!���,<4�9>F���&s��9__�4Z�����ώ�2�iR��w���, ���Q]/U{�b��9XеțNm��2�K����߯��[����i���מi�ښ�2�!�fM�va�;��>��,a&���E��ub,���q��Ed��\�+�Aw���x~��J=������h�l�V��$a��=`�nL�$O>>��*��,̪l��{P�}t��^���=��X�i�� �,�n@��c�N��W�_�4���B`R5�U��3.��~XւT� ̌U���t?��Ih���~�=B8e�2���C�W�EՅ�
HH+H3HwH7"� ) ݝ� 50� �4(���tw
Hw5 ]���gx��;��Ώ�����{�ZϺ�������#�@�Y}p����s���RI�w�3HR�(=�v�m"ׄ�r]� u(|�����7���o�;����ݚ'͚վ}~�=@�_}�1��.R�ƹ1�m�y_���(�O��-N�/�j$�{o��7^gdg%g��m͍��������ر:6�V�v��"E0��]������R���m�$S���x����7���6#.��XX�g���M���%�}�}2Ԋ�>�#��L�ч��a���n�7w[gw���U�J��}r:YH�"�K�;�OSs/BZ~�����K|��l�����S1(��8���d�ӊ���5q��&(5�{T���)+g�I�2	I=w���7 �
ny�!7~��E�P��+o ��ݧ��|9���#���"��1zO5��u�����u�fϒ_Э�$k�zL̓[9�q��
It���֙�˭��Z%�`>�Nm�N��U�,�R�� +/X:�#)N��UK���C1��|{��|���`QzŚ������J�*�&�dƠ3RN��^���i��뀼LsX�5�㴬�j�BX�LRr~a����?P꩔�8(��d	��1s�Ȅ��yor�.Q,ɶ�<e���o����Q��0��6Zf׌}B�}��⚱~��v���o���'�A
�3f�N54�_��0�l�k�_=vx�(�TB�%&`�����B��1o�;�D�G���e嗙��A��1��E���߆]��s��P	m2*I���9-�G}���9����_ٌ��:��@���߮�w�gM�*��d���^:�b��{�AZ��8˝O�-�Q
��������, �9{�Al�h+�M���g��,���
.I�(ӳ�.��6���/�`ϐ�]1\X$������`fD�w���
8�d��5zG!��d��m+>�	|�xu�U��D=���6�m�`��;������������e���Ý�U7�����u*���L�|TC�?\�*�13�d��K���~4c�c(/��hP�i]��'��;��0���lK���h�=��E�[���6�߆��&�Ř�g�$�w��D��3�YU ���J����U�&/L������+L����Ò��r?�����a�^�����$&[M�+�����x@�x&���ч�|��,�mt�6�^&&��,���y�9t�)��3=I;wcmɻ�y>,�W�(�����n��W�\;6)-���RhħZ�F�M��P������}bq�YWD�����@G>�Z�:>��ԷO��q2����&�V��އ[;q�j�|��?WT5I�8LNB���D�?�j�u~V�.^�HuI�q�҇�vM���{���$K�P�?�/�R�f:�����ؖs�P�ޅ�6SH�=���=�Q���(�*O�2ҳ�+�������Vm�� [�$
j��r����^��%_���\�A\H�h0C�@oK	N|����޲�1�+��\�Z�$�5���y��{�HuS�Z�N��ڈ������0��fZ�GD��ZF�=����tk(��ѕ"Q=�Yi��w���M䌰;�-�����ـ��<�2 ��U���|w�<o��j�K������v�oY�)/?��#�;��'�B�|��~���ݲ?,��D�+�O�\�b�g�ݜ������VWF;KvP2�{Ղνy�QQ�!J,�/$���ڛ��LǏ>!I]B���W���aUBL�ʶ?Hr�^��{ؤa7G�s}���01�������wiOHI�Z�i;����.2,�5���2�`>��n��S\�P@L�o��1�t���'�?|���t-��L$��Ck$�[D�r٨�w�#bU��]��;��͵ܮ�_%�0=�N��~Z`�!�h�����ƻ#3��D�gXf�����~F��YZ<���ϗ:��c��տ.��7���)/-�!��h-��6�������ZZ�iZ�"���ʕ�R4R�f��|#+�֨x(��L�k*0��Λ�T�,�m�$e�C�Bc�k�e`"��@�P}2o���5B�=���5|4C��a�}K��yu_+e4_Ë$
�,�B�f4�x/�&����k�0,������/� *Q6� ok�vqw�L�f/��� [�l@s�;�j�n׾�t��3���WO\8?�΅�x�6�,��D���c�#n�6Z��ssiדN�e۲D�lr]�2�Sn�a���W�+K�[��U��8|� ��W�4�!Z��r�K�F��b��x=���v��\�����4V��'Ը��uw[�T��G \b̟��8xK"��zN�)g}#���1H�3����a|~
�L�h5j�D~���O�S-�3vy�]#�?��8���"f�����ڂ����KWM���S��%������]*�Z�j���G�J�J���?��,���[9�A����Qţ6P'����yB�OQ�yOt��[�V]��kEG�Ŷ�AM���7�+lƈj]���"�1[���v��Ҹ��ޏ�P;zf��6�`�W�$�\Yo�dt
��y�>엛�ټg���=^h�瞐�b*������D���/X�dݠ�r!ԩ ���$E;N�,�s|�j%L�L�D�����w�?ih�ҳ�_�r.�]̬?���{L�� Ӿ��ǖ�й�ډ5|�����a���Gt�S'F��i��OК�93�d ��Yö�Ǧ�l�=_��x,��#���鸀��w�Ѭ1G�nо���+3.��u�ɏ[��?0h47g|2E�f�	F���Ȉwu8|�H�5-P(*�Z�l#�:`;- �!��򥬶T�rkaώ\Oia���^�W���Ԕfb'�����-�Jn{��;ӱ�cG�;���0~�L�lcF�k��⢗��
|�V�� ��s����V�)��`>�Jsi�ZZ�1ɾ��3�e���x��Ew0��s���JN�Ǡ�%��AU�ٱ��= T���"� ���!>���ٞ����S`�_�'4F����D�������}�rۭ��!�~G���<�z3�{���?��`��;��9jsW_w��6Ȉ�w��a��yY/�2����,���[n��"��"��͘{��҅
�R�螃2q���w$>���#�C�M�Vx�����;�ѕ"��ryz�`\�����?d�L�4�2�zd��v!��tpEǪ2��8`�3|?��Ԟ�ǡ�1Z�E���Ul?Gt6On{9�!J&GS�L�G��KK�!ߗ�`��s��K�:�&�9�@:�l�i"	�8��ذ�����4�D�r��CHs(6d��^���}̕a�l8|������[�P"�(�q��㗯��:T/ڂ��=��4]VF�� l�;f����τ�!$L?+��N��'�aH��>���'����dIZd����ņ���F���YsH[�i/�M��;oy�۞���豶�ű���'+��v�D�X8�D�z����#��ί�N}b��L.�L�	u��OK�dJ�}�����R-=&�����73�f�a�]O�6�\HNLׯH��n���x�m��Ș�d*_�c����?���b���75����R��ᶎ�Hc�28�=�Clef1�ǰ�򥸬@_t�@���5PX�Y��h�L�/���f�v�~�����D����5�3|C:bz�5��v����=M:���EM��ƗX��5�,M�O��Q��;�O��=Pp;�Dc�O��(B�Z ؒ�ʆ_֗����9����zF�3C���cZ3��U"��FA����E��R�%We7 ��'L��ń�_pb=������Q�ur���w�"��g��=�[�|�� &^A1f���0�p�E�����y�a��C"������J�> f!��Dc���*mܥ���Z̪�0�,��R�o�1s<mk#ZX�:���u��/*��j�u�K�t1��h}�O�jZ��̷G�@g������=���=D��8��%���`�ʶ	������i�z�iu]V� ��do��)���q�.�/R~h� �k��ƤX���kM�?�o��Ho&˗���!g�70����#k/��H��&|��*x'(���Ѽ�����p��I�E�"��,MRl�d��]Iu�7�'^��T/�kg�ś� �-|��:��>�!���EyR���1Z޵B��P蠮\�)�@���Ҝ� ��%���p�M��4�|��
��2ʚX�,�4��Ql/eQ۾i�;�UDu�h����y����[{;��\ss ~��dR�����{��L�T����H��z��Su������c]
�ёjIޚ�p�:���5��[%r�0[
��l��@�q�k�6��C��pM�/ɻ[��yl��1ĕ3����:0�R��AsVڸ��w�����ɑ)o�T�E�,>F�<$�ѷ3*��f��|�]�	��@(��z ��\:$��E5p���\0��S�_yY%��*"���=��;��(4~8:fB�]�{?۾�+ OoR��' �� ��d����[jZ5�i������VԦ�l���w���(N��������Q�AO��f�)��Y�Y�����=� �����`������[��m�-�ӵ���ѩ#���/�#�It拼5!�Dc	i��Q�� B]�����e�?	�@��! ��ó���6�-
���-�f�컝� 2L��z2c��:�X���ɔ̈́��}�KA��[��x�i�{�Rq�A��F�N&,3�وj��TM���fbZ�t�Ǝ:K�^C~o/6�f+N�����7�ui�I6rq�nR</�P��!����O!۹	�l�۴2Ap�p>s�û������e�>Y۱�d|���իB�`}�R��c9�腩G���?~��?^�z���p]$o��!�w��;9�y�)KE����bY&�ػB0��ه�����j���,n�Յq���Οd�pP����iT۵��9ڄz1�P���MǊY=%ТL�}c/���F3�_�sJ6��9<�����s��U�����kqy��n�+�p\���j}aLi�>�q���0�n?`~7y���w�g4@&?�)����<������U(~l8�o��nXY[���X�"Z�ۀ��ܩ�e��H�a�y(����Ǉ3���C
]��5Ry\��œ-�-X�YdU��zq���pܔ=����iH��Q>l��M޿�C=���tn̢�n��?�B���=���&/o�i����H~]'W�e���EZ_F�F�Ё�9�Ȥ�g:-wOf�gWs�Q����2��'�%|�,������Nkmɠ���em�/g�������Ԇ[{�-N�6���k��l�a-˹v6ij�w/80��4�ND��������oaL؃eZ�#B�/:ߦ�ކ��i�*��^�l����塞�����q=���l�.�V�x�B!IR���2/���V���&_P�ڵn϶����0�6���ٜ�����xB粔�`�~��%�nIA����Z���ܥb����1�Wd!h����ف�%��e��{�UϙNWs��)-l�9S�k�����o�������­����|b��Y����'m��1w�w���,'W�)i���ʵ�������q"��H,�נ�����B�<k(Dҍ:l�U���ˏ�{J���k>ď�,*��Ɓ��!+��p	�/Gq`d3����������,�����>s9g�jhn˥a�!��aITTZ�����x����\BǙ铿q�m�vT�O�B�?�d$P�����N�_l��{C?�!���TWc���+zs��P?m�#~��wK�હ���P���#�Go�lR�&�>�ۢHzQ	e�oH���wT?>���OLL��!�OxJwPE�]D��i�x�M���܇"��@����>RF{�3��Jˑ��C֛���S�0Fr<���$g�?`�B+	w"����Iiw�m
s	anr�����5�_�� ���(��/��9��\�l�s(��y���=/�n����x��h�7G��߈=t3����|t=B�w�J�ujʹ �����g��h
��ٜ�^k
���hE�U9���>H���糭��tr����KC�i���{��>��<!�#Ak�ӏ
cIF����sܕ K΢��ٝ����lO�$���R|��/�=�Q�;���~�i���1z�����bzz3�Fo�0���}�Н��b����BS�%������4�:XLU����ji�x"N��o�;����^��5Y*�k�)������M��#�vFY\?-WaU�OQ	t����nY��Fvb_ފ}~����ZMW!xe�r-|�.y�r/2N<�p�y�}d�I����_�2��a$�N'V/7`6q��M�O�0� ��e>������.���vEW��_�wpq�ōe�U��v�^{�hrt%t�6�ps�"M���C�3�t�d�?��� ����zJ���S��CZ�K����f���{�m��b��Ό���+������h|�hf ��QES�f��nH���M�D(j��e2��R�Cl�-W��D����[.���0��d*��f�p0z�d�������rX�Y ���N�N������g����J +�|(zB�=��Z �]�!�pèn�V��Z�֪�J��=A�����S!�+��)N��:����ċ���cK�7g�Q9�[0�+g�mo4���2'���cZ[%l�=�!�������(�P�ۜ:�xO�V$��,G�$z3z`�)n����J��TJ�}-��x�*��1��B.S��{U,T?dO&!��cb��]��!,�uns�c�7�TK���7uFY,˄j�z�yF�Ɋ��)�gy���t(2�F��ǔ�!
�_��̪�'�_�8����8�4�������ߍ�n��T��z��EGO����M2��U��,&$\W��/����6P�X2/W��kQ�,��Nq 6�0�kЃj���i����/��[���v�.$���W8�D*��u(��?~H�F9κ��E��T�JЙ�=�7wy1ə�2��n�d� Hu���sZ��B�GQ�;��z��!B.�T���{�,g�e���Ч����n�99:F�IagD1>d��ˍ��n�vV�{V���HC�����qe���J`-�f�kWP�M���;��/��!���7kMs�
�'��k���{�����+t{t�W��W�u���]��Ŷ��
��������$��C�a�X�B�:}��]�����Y(y8c`�|� ���%8��%�X#�^02�Tl5�JN��r�2�tf��re���X�ߜ�#�!ӣ���W��Ch#�'�_��A1֑�(��B����ﭽk�I����K���:1�����Z�K;�����e+p.a��]	<�%V����5����Wk�LJ�G��_�^r�l��~��k�̙�dc��
��u�'��4��";ۧ�mz����oQ�՞�����/������?>A�fr��}���~�%G��2��hA����)�1�T�u����:�h��2�+g�v(�X\\m�_�j) F̏��r�M&������0@�*vʇ'�{J1���Y/�D�+�q��r�LA�h��Ͱ�2
����K��%^����*Y� �RMq��jԀ�[/bFz�r�Y��^�������v�����v�ڻ��5a'S����|����ؖO\|����b�7�Ga�d
���1ؗ��=����<RX[��Y��U�B�8R	Gl���$���l��j��� �b����UV��aW]��͞��Q����I��MR5���LL_l��e;r�?�5E�*,���Y�Ƕ��������|H�t!55_yƆ>S�`[���Կٽ��o�~�-D�&�O#2�W�Qz%�����v;H���
|�y"޵sap;�&��;��#3�\��\�U�w��[e���������*-&���V�sn��~���j�Ů����<Mf�o������1�.7�o�k^az�+���5�n���"6�7���}�n����!�3��^�s^n#�ۭү�FN����'��dJ~\/�<J�(El��*/�\�^YJ����TY��MU[r)k���O�?�V'zw�Ip_�ح�3�c�/���i�1gl0�a�V�Pl{vd��DP�/-.G0!ևpG�cX%tl$t�ȇ�7�Zv�����+)�����v-N+}�a -G�l�Q��s��=��C(r���u�1�,h pW��z*�����2q侢Nk�클�|��$�FT٠:c�ҡK�U%�%0u�J�h����u�G�0Q�<�J.Q��I�F,|I�`+�/���#20�磷Ѐ�g�	���ƕr�;9�F��E����wY�VY��}	jXi��A<�uu&���b��3���J�^)3y{�6���3o8{�����rf�9�t� MR>PW�]��?[;�Y�S�'jˈ���9�!�9	b���p�p#r�:?55���o%>��UL.I�|�ٌ���dEbn"7a����}�� ���:�:;|a�a�$�Y���"�z�ؐ%�hW(w_a�Ylp� �\���Lx1=�,�h��雍�{ל�ސ&�e��?�BC�M5U$��D01PPܞs^Ѯ��?�+"�!�.��p��Ni������5|��f�B7��\�h�v.Ӕ8�&H�|c!���&�%�GՑ�d�#�09��5�O�GR�{��&�>@����`3{�t�?A�=9G��~�3X����8pF���w��6Cn ����EH�>H�Ŷߣb��P�F�x����kv}�G�����'3?%6��R�r;�dv����
L�Y�ilȃ��r"o�_�-D`��v��<��7&�|l?�#�y"�-�n�����wT}%,��a�!�&l`v.�����Ix�>"^��j���	�\���C�I���y�v��6�DEK}�#r0�7����"P��k)n>cU�`�Zn%񂍰t)��	]�L�2_�ݭO�s�r�-�elM��3�g��û�-�� ɧ#�c���������Eɼ�eJ��B�!�]T_����<�z�T�9��k�J��~N|�e���B�=tkF�B}u�9NL�W�ҽ+ة�{��	"iugt��޿[9�<h|a�"�=v�z^eE=xS��9K�6�TL��}����B�tek��h��Mm�S3쮸����r �������K�8�O�D�����Ѩ�[0l������ȑmؐ�����B`ɀ�3;oՎ������$6��Q7<��\�ܲ�9-!c,m��A���$]��a�y��N���Q�� ��#�>G�Z��� �y��d4���CP���PevZ���(j��,4=7���ZVfF�|/�����#�!g�o�є�"핌9����z�`�c/�n�U�"��r��l{ȁ�A��%����'{g�%��ʑ9���s����ںWG"��h�1��A���2�A�A���sB�`�J��g���D/�oŜ��1X�������B�1r�\�˯�h��Z�ס����������7����w��I�&��TBVVT�>�<a��3��:�\(��6��=]� �!�y �� 7��)���fQ@`�Ҍ{��>@a���˴@�K�D/���KK����*i��ݬ�E�ڴ���#g�!zIP�aϳ8�^��j�#��g	�7��f��ŰQ�Z�7��1����'U������^^f��V�����Gq�Q�X�u�Q~�~;yLt�g�!�`���b;m�}P]/�<�PP����~�k^ ZM�j�^�KK5�a4�acA@�qP
�X?�7�h.&V�w��b7�ӽj�SY:g�R5枉a�V�<Tc��E{��!�z���l�8	?�����_a=��/�l[ё�O��j��G�P����om/ץ��˯Fs���i`��g-�%��ۃ�S�▯��R����pH|-ǖ��\{ ]��(@~E��j~�������Pr�Կ�H^��fB�cA._�Ӆ^X��HN��]��W��n�$���F{nd%�54UX!�k ��Xq
�j���w*ʻ��������e�j<���?
#�+V�ƙ�t��iP�>Է�p*\(g�c�|���z+�{X��)8R��$_A�]�Z��M�P�j�"��7�uIJ nسna��j���Pd���an��`��cv��Z0x�V�Z%��A�9�o��׊h�"�Ȼ�$�_t��}������>|���w�݋f����g�����e5��Vñ;�~[g�CE_��:���&�wm�S}n������8Z�?�K7q�>��Zfk,��vh���}�5pF�7��p;�c�^��[hx&���k���!��ro(��;{���׽�d�)��O����#�k�2�	a
ڑY�ޭw2�* �Q���B#7�V9�x�s�R�8�����'���&�/�-�@���
�[N�� .U�+��݂��Rrn�����+��ؓQ�`[҈���#��!G����/��^����դ *�W[[h�����hR�s�Ȅ���pv����S� 1�#��y���34]�P�b��ͺU��~�B���C�������ɳ�7�:j��g;���k.=a���������v��ސd��#	z�L���"o��c�]S��h^.W�d��#�~U�˴6�-�KIO�	ށ����d=d�[��Nː�y��a�B�����i���]��\[nN9��6�/��-�D9�������=�k����W\C�`�WX2d)��,J���Ei��ڠ@'P��84Qx�v�6}��-<Cz?�彧�.��a .�a��v�?%Fx���|�����^.��W^�������X%u���uZ�p�'�9�0�J�s���4�~�t��=2�����5Gv�X��e���eW/�T�=���E��Y����䵮^��R~o4��28ͩݚ���uZ.R@�w�K��� �D�����1,��U�iy�e>eY���%��K+Z�4L|@�Ob��&Yc��h�M��uD�mjm����-�q={�)3w��C���Ú���8�:���JV_R2�q]F?92M�6�������(,"�ϋ�T�Υ�9rz���g�3ҹ�K������ٳz�Q��ښ��a�ּ]���ޣE�&QC���"c�1=0�T����w��m��Z?�i�NO����T��*V��(܋��,DFIw�*��O�3MA�8�U|���t��
D��n�������,B�t��d�E�1�\~Qat� oHh
�����Gd�c��P�Y3� �>�Ȕ�$���������˥�q{��������cfXM'�0&�]�d�z��O�6�r�"d�%,2�}>������B��Ǣk9"���2g�k��C4���m�AK��""P�-,�-f��}�fR= �غ�;�ȴ#�r���࢞�ޜ�q� �A0����]|���r��!��mU���+؏|^ɋ�/��̟�/���^�-��DB���u�aE�:
H#_E4C? 5C���[�a՘Q�[Q8E��Ԭu}I���X�[�J%�N�ȵM�Vh�>�K����M�/'dΗ������X���e)8�ɍ�&���0-�O@K�C�� ~�Z����p��������uz`����������^6����I�ä=<���n��Z��H��`!�_�Y��M��
@������:K(XD�cNB4u ��Im���¨SpS�����2�)�|<��!n���RBC��$m<z�F)}���c�7N�4�iW������Z�|�x���k'�a��b�{(Ի >(a9��S����PmѢ���1i���veҲv���ZRg� d�3�C>� ~�[R��ș�-�sh����F��Վ�wC�eX����Z�$m*@�](QO����G�)Q�s�B�_�icy��%��+���l,����E[%�������|�0�$zj�Y�G��E�(Q9'���:Io>�l@$�Vw�)y`~�$�����	���ǿy�Et�<g ����/���yhVu(�b�����,��Q#�h�D�I����R7xՙ%-:^�ƨ�T>I�oh+���/�,P&�$�o"O����[��'�	#x���)QZ��T����U�����]�'r䜐qx�g����������g�uOɴn���U4ղ�ag�W>Y�-�a��X
&���T�z���+Mb�6��̬�V�'��(�2�>�_�3��:l�RM�#^)##�G��{�J���[���ԃPP%-e��<�;�[o���;�jc���Z����ϕ�ȷ�X58�h]�z��=$��{0��=�\����F���ׇ����&�)ç
Esn��t%ݝ(��|Q��1m~Ǔ^|"��I7��&ܘ��ؗ-\#ddO�=��L�܃��?%��]�����e`���ƟW�ܠ�@���%Ep�OD��`WL���*�q��t�,B������e�X��yS��Q#�en����ֿ�4��9/,y�F>l�&#K������Ӄ���Ȏ���a�Vo����t<��h����0���rK����}׻:�����E��"�(S�EI�C��;V<C��Q����CO\267�Yqpt�� �VP�'k��'�LAf��,��D]v���+�?�����9��g��*=�d�03�8p�/UbY�L�Cq?Μ�����Wh~��uH�	}�b�! ��bD{ÃҚC;hy:qqy\E�`��A�v&��{�0hD;�b�<�]���[��v��􌈞�q���.�Nv��R�8���fZхQ�ߓ���ݦ�1�	�9ы�s.��]G�����t�u����4q�
�~�5
�0�$��vM��g����i|(3-���'�A��3�B{�O�D�^�f���Mo�!�S�䐺¯m�ˑ�<�2�AsK�<���t�F�Fe��]p�()�3�k��y�Ϣ�Q
!���Fyf�={�eZ���5�jϣ�W�k]6��J���w�(�ߺ�o�$U5���=7���ǫ<@he�\�)���;�����s�p�.!�Q�}/���X���a�Փr���_�b�$�6���Nx6�e����U��3���Hi���̶]g}�A'�������1�.P������c�%���yg���A�>�6������~�MO�&��mJM�d��ZZ�gW~�b����Gy+\i>���◎%��������y�Ͳh{�}	W�&�,FMlM�}�A��2�<��Ũ� �3Cz*��'=����,�-�8���R@�N4��Y65Y�`���DWfڔ���Q��Ȗ*S
�	�<@�vw���� ��ꩪ����pa8߼���Q�\ШS�_��dl�GO�w��ݪȒ~�N�PAL����&E`g�
��#�����%f�Ъ�.�~��T9����7�
����ǈ�^��]��e͟/��\�jgh�7�N��"�U� ��8ʀE�L����:�����?�����þ�.aŘe5��
ｭ ����`���&��l�5}�7����7�����FS�@c��|��I�h$c��d6��9����{�RM��������1�No��*v�FL����I�&XT��} ɠ���+��P��#$��o���TjR��rs1^Z�v�p��`T9(h��LUg{�f�!i|s�I��`���HYh����jA��k���"�w.Vf,�U3E3�����y�t��/���D�k,�d67��Fv_ҿ5�r��]�Q���C���ZNo7,E���{�[����8�5w�ޫ�C�a�!��Ez�*�5G�^]JĦ����e`3L��ʱ`!�r?�e���L��/���Pl�68���8l�%q������(9�v2�R}���u�����W����FT��<�L�\���f���(+��x��K�y��(c6�9�]mg/ӿ����+"��Q�m�D�;9(��q����dn�!ֺ��+��/^yUː�nVd~v�t0T�6r]p?�nQ^Go��b�7Ҩ�=�Y��u��|y��AKG��n����>��]�������/�2���1�| �h��]�yr����5O��Ts�L �M*���&c��Xl�
�1��o�޽0e����(k;.�H]��2Ly�fն�X��$=��?>{U�&@Y=�;�<����g��o����B�^BJ��0�r��B�C�����.�Tߞ�tT:�lL&�"���9O/;�d:�������k?q����.�U>y݁���{�K'�U���PN ���=�~�,**F�pg��������מ��l:kB:����)[ܭ�E�糭��+�+��G)���r}%S�'ss?3�T̊�����˪�}����Lo��b����]���]N�_B�|jo1�^�}v\��}�WZX!ՒQ�(��;K ?�G�G�C��/e��9����Ol�a<h'A�a�����g��������n����݆�g���g�_��u��������SխC�C���q\WM��2y��,Ug)MЃ���@��o�wjF����\�M��jE�9-y��mM�?�O���gGh��j���yB���.��Ҕ���6�|�_�,�$eeu���9�W�9��)�{�ݻ"�ϟ#��E:$�~޽:�;|{�0�.�� �@�(�s�4��*�����oJ��5@��U���RX@ߺ^�/�*�A��/����"g�[J��~�j՟�}��."�o�z��H�#�?n�⾑�Qu��h9Ӕ?-֚�^b�������S$�k�vY�9�O�U7M�м�%K����&��y��in�ز+X�hw����}�?���ccc�.�dP猾k�T���Q4�ٳ���V��kP>���x���u�:�Ўh��o�f|�N��7�C46�',56��7��.����c�*;CE�����F����#W��~ǃ;2c�v$ʰ�����z�iͮ�E�Jq,Wb��-drX�7ғ�1SO��X��>��������[�v�{�8�wBD����ث����~��Q<�-�XnYk{�:��n��~���W��Y�=y���?���	c[�J8���1�g��;ei�� ӆ�Ag����C��b���	� �?!
��5�a��ї�#$�O�xI���~o�PR�̩�BIM)�аFc�ι�� �X#X����ׇ�8�D4� i�:�(e�ϱk����4	�F C�E�~z��D��M$'H��3���oyDA�P�as���U���a�$��o�#�s�3��$-�A�s��ߪ�gG��"̞��:o�'nT#F�������ܥ�l֏��f���/�JS(�$�Z;R��Y󄑎��\�!~r�#,kT7L t�殮E:e]�@�/�ԧB�F?��+n/d��ɺ{pP'~(״	�AǮ�
E�?��K[�`��l��p�AF2��R�#9l$��-!�N��ߤ�a���n�����x����&ٮ��p��Û���9&S����k�{p輳��R`D��cWx" k��s��-����\��U���%�q�+v�o �8����-���u[���7����Ͳ+UQX��`꼅A>�Z�.����mc|�WlT`���l�H��H}5]뢖���R"=�r�c��(�����@#t����m��47]k�zR5C���o��mwL�lK�`	f��X|líH}�^�:�1`�'�$�c��������-D�'��C)[Q��g�Ԃ��o��͵_�����-n ��q#����ݵ�s��e�De�+$m�25#��.�X]�ZY_�3�a �g�,L��z�i��%1�����=k�feЙi+��_%���>�>ҩic�����T}K��_��m�f����9���󣘨�d-�n,��AZ���Ã�7E�u״1y['e�QM E2�3��5�N�ըV_�Oװ�6��N�HVww{����Z��ڞ����F;�3i�����3��
fS�n��Ӿ�P�Yw�0�R��_ش�tew��k&���#����.߈�_�[]����mMèN�(>G��3b���h���i=g��o~kB��6�P�����r��no}I?�<�gQ(��\^-H��`$�Ԁ=��)�^��%�b�~��|�#��K�~ϒ�Y�J�R�����)�%�沴 n�((��;J��:�i�9�����.����;�	�F@�l��B���`/c��;RY8K�DT�ur�v��8��E�
)9�aX�:��gFu~0~ �΢T�c��d[�f����^H��&ge����X����/���'�����mW�o
�:���Z���S��G���J�\�3��\�����0�VF���5��� ƗO��:RU��R�>ܫa�Ϻ��ߟ��������>�qS!�D�7�W��|�a Y����X��`�\�TU+0'��:$��f43������.H��4G�V�M��ʯ�bo�&Q*a`*t�8sB�)��^��=��t"�َ��g\XSN/�6XD&�Z�ݹ�����Y�����'�ue�!�u���F�,n;��������Da� `��6 K�\P��������� A �������V�rM�G�����c_'$^�����
;�Xn� �ݬ0���03$/�U� �Ŗ��kq�1i��ڸ�6[����^7А��N��\���FN��'9Y�Q��j�]X'����[�4��B ��=w.��Cpwww�=��N�;,����-�,,�G��w����ڪݪ����9}�LWw��Y���H� }w
���� r�6Y��!z��!k?�O�0��mX?>X��0@��M�L2ߡ�wd�o&�<���i b��L��ϗ��^�ʽ��y#^(�����}��q�q~��`Λ�#ֳ��_������T�u�+�rk����g�����u�J��Ï����h�k1�{i9� K��G��������PX��N��	�X=?�����V�Ջ(J�ԛH(�%S�?,��J��I��+���h�tw��F�� �i�J��ZoqbbAkc.���և��Q���w�~6��7��r9���[�l6��vt�'���|�PϏ�e$ZZ�(�P3��(`��X��[� ��'{ 6҄
�o>
��SK��*����r:B*�y.����u+]�p������ZqԗS���TRV����
�wW��Xb]�z�;ק]�f�lo'�G�vQe�_[���.ڞ3��[yxҼ���)EW�Ŕ��.�� ȃ��,��R��O�ö�ML��%s2`^�H"��~�%����+�sӮl!�������������E�Y��⃃̀:��䬯 �R�X~��"�O���	�[8ik{;w�nM�
�겞qs��o���0��jꓽ~���xjz��ื~���f/�J��x��q�g3���3�jAE��ײb�ӹ'�\��)�+x"˼�@�}��qnJ��vL���#mt=���g���q�$�����6�GNʸ�5���������nD֙���c։v�����K�0Bu��س�DǢ��a�X��_�_��(n�����OC�9ҞHՏx�R����=\�����x.��T62�Xm:� ���5�Ch��f��N����%�;���w5�}�P^O����O�&�y��~���:�@�.�Y8����\
���gi��D�xҔ��nz�t�^#8�t��f<;�vh
ߘ����G�kQ
Ú�F�rb�4-�C��T����9T	sUQ(���>�͡���x��qy�8�.x�|\���7s�7':��6�c�@�j+�������4���y+����͢u�������H��Ϲ����G��km�hXΡb�A�q�!���Q���E4>�n��!�üj5��3�@�n��5�46 �8��;�fKC�W�e_'ؚ��F_�-x���m��(6ā����<��ǘ��&'qu]��	��Sc;�����|/5������΁5Di#}�b 6���L��;���ɴ�w���B�oYO��e5׼���Z��nbdU�U���3�]�T�p�T�G���h���Ĝ���Y)a(��>����}I&'iI���l���j�	���%�+y(?K��'%f-�iꛤ|>���3'��E�*��&7܁ 0��/;]kum,c!-V����sނL�0���"����XD��/��)Ö8��m�0y�ԂN��J�'�y�*�9�-��Fٹ^ߵ,I(���І�^+Nl����F��q�o�:�Ǒ9i�i	��y������v��dy���C�Emf��tLm� Ȯ�����+(�ݞ=}W��J�z��|�F���k�6����!_;�K�x�R���8��c9����_���(���HC4#Nk$�.�P5փ슓@O�����e�b�]��[��k�b;�LjW�EE]o	Y	���wmy\�c���hq���à]
+� e��3�ς:��V�՞�8}EOꮭ��1�-��c�)#>Ŗ�;9��_�4~C4r�{�!;�-%Y�d&:����7�7GYv��#��@�x���JԞf�t�16� �ם�u���(g���ŏ<�p���6�Ԭ�u�V�l|�m�BD��h������BY T�	ر&�w~p�c���&���/�1��yr�1��L��'�]w����I2�������F����<}��8�y|����)��	̐�q׾�潡�4�0pw����xQ݀sR,O�h�dzy|��׍}��^�1d���M�;�E��g5� ��h@��CLe��� ������'�V�2�LF�ye7	m��f"º�y\���ǂ�$#Ŕ�i�#�Q�g�c�7�����Db�z,S�}Ŏ�UW�-��(E2ooG���0c�J���4e%��/o.�}(6�Pd�-4C�r���y�=�'��͒�k�IY�?EIz�^��O������D��><D
RWQ�c��	�Π�j:g.$�l|[�}6�Ϫ��J,�.�<
����]1�*�U���Y��S)�(�&
c��5�c�N*Κ,P�H@������p��s���/��d�@sT����M\���/��V~/;��觼�E�V�0;RKu�\!D$��M�w?%��M��/-�w�}�޳�R
����3��ѱ�^�qU����| 7%�
'.='�/���i�`�^�A�9!4�4�K��X�du�;���a���E�Z��{�w�&����~��X���2�6#���O��5E.O6�r�r�aIщN�i�|�h�)R,��W;�mv/O��Jd2[��NHl�+�c
I��:��C��?���ϺmKi  lq\���G�R��9r��b %��E��F�Nx�uq�E�H0�x������2V��v���2�� 9Gv�O2AK���mjJ�M?W���R rƒP�V��("�J���1�,4�������~�T�����~A"��m�;�;ߩ~��a^X-REa�m��)��r�5#�ksyK��Z:�JM6�l��w9g1�o�֬+�_����|Pd/ɇS'ޅX�y���a�DX<����z�� ��舴�dsL�N�n�[h9K�qh{��7�K���[���	�u� ��=m�4�rVݾ���@�U��
�7��-�ى����㋊&ap���[Gm��;���؇��*��i)�`�cpo4�H��?oFq��Vmпn����x�c�״A��ė��㰛�F|M� �z�=xCL���O�+�U�n�v������K����j��F���sjL�p�g�+L���%���Rl�f�������h��I���/y���F�E��K]�A�>��h*�4G�x��LL�5���؞-��c�3��u�Q�V���*���#���)?R�~����;NG<J��kp�0u{W�H��'[�C�� �b_5i�Wy:�)=�_r�L���e[;bE���>��J�oIoz�ə-��_X�CR�_��we�G�'�Ob)�������/!��b~x ͧ���x:F���b�Ԋ%��OI��Dee�{��U����� ���z�g�R�>ɊCq	����٧^Â
D�}N��t� ���U?���B�5ỹ?�ج�V�,W�W<�Y��ݹV�O�?��8{Js2МG��	ox]�(�Z�g+��x���#
����ԗ�`�Y��������i�#�+�e+}1���{m �++<R�xK2�&���Sl���J�k��۶ۀ�?R���R���8R�-PTjUq��C����L�����m�-[lS����n��bԩ�n�"u�>�7*W/5]������}�O�g����'c&/���� �,��7�w��&8C�3�W�2������\�D�Z�Ǭ;� �w:!A���H)"��k��ǁX�N��B�|jhq��*��I�(��#�
E��^���o���p�U_Ojի�5�}�nM����g��N��v���l��ƙ�n��أU�}�b���6���[��ޏ���h�*�����0�����X�l�V�+\�2�������url�kD*��p��a�Gf8�Sd�ek��V�:����PQ,��"8I�jWR�9�/���o̃�.h����	a�D��#�E����}�u�l�&�ﯺ��lh�Z9�kf�K�R!��nf �I��=��|��A�r�s�hI'�������Zg��`�D�JG���3ܚ˩_���-A���%�n��wE�t�!���Daձq}�!*��J��m�
9�����M�R�l��ť��U`ÕW�~�����@��;���a��n
��l�j�x�p��;���2��T���,�Z��$Q+�F}4KSUd�3�-�i����@a�ѳ'����P�'���;�X�+��^c�n,āNP4ㄘΝ�<�0�My�Z�s�%s	�[��frq6v��D�����[.	��j��˒�>�J���t��w;��.��N�e�nZ5Y9�(s^�����d�/�e��L�:e�|N���#�d5�:aC΅�;�2�����?����,�yOh��o����|=j���|GL?�ߜ��� �(�V�g�2�׵����Ǔ��H�>G:�Ulhv�bg�2z��&�LtӉ�AV|4��t� ���z[��ܔE7,�2�y*��͞2�9^(D�[��uq�/9w7i��]HOgF�i��q!η<��չl�a3
�ȵk�:��Ңq-}�+�	�u3�Ӿ��y����0>+�"��D�E�U�`,��nlc+���"mj ��Ū?\�.�M�^�?���Zܘ��nd�6X �A5�3E���l�v�P��}�y���s�yg�)S��|�stg� ��/W���pq=M�Ⅺ@P��o�u<s�F>�c������_�]##�Zn3��g��?�����c�s�#�e�K�[z���fUE�S�3���$P5}E"��z=�p�_qh�&Ƴ�S���i�P�\�ݥ,>u)�b��;C�eH�@�*B��V��(�Q�Wnf�R�~������+>2��D�/���"���t�p�{a��,�Ĭ&�L1��W�-^J?Ӎ�L��5M�	/���V��8}�&OA��f�ɉe��M�U`��,�O����B�����֥P76��4��i+�:����am}�N�?E��� �����B�0X�K6og"���~�	�!�ݜ��'��r�9���PF
]�+���͝�m���GR�7��wQ�bog2�b�n6����%�P��#�?��Z��I�ys��Rf�bOO"��ʲ~xa�����X0�o����n��"�
G�v�z����+b�{�K���Ո"{]�CF+k�*�z�kTɛ��)"bl3�+.��[�;�AP",J;+�4�?�x'�[j��G�"��o�%��Q�p�5q��>p�rO��v�T]���u�@(��K�V_��vۼ�_-�9����c3�j��>!1�㪃+&I�Y�Z�n����v����3���ى xu��切�6���{͗��|߱�V q�����}�BEXi��Z��lf��a�jT��{����;e+�2b��(���Q��%�|���@�p^mՙ�<����="���*g�>�W�6�����%�`�ȉ�ޚ��/:��<s=��c��f�hC�jF���>ߌ��A������߮�TE�b��1��؄�Ş�ܺ{���)ۊ���[ƶ��S<~�ޟ�( �.ip�����	�4DSX�Um���q��i4�P��A2��.��S��/9.�����0�h!��.�~,�In�;��)f������m�p����U�|l"h�U��^ �Խ�f[��ڛ:~=��B:��ۚ�����D�Ѹtd�ػ���Z��������ƞ��𩯖�߻��-�Z���
rlq���"CN����8�Օ�|P�o;�v��C�_�����<���UU����٩�J�,��X��̴#v�L��b���־�P����Sj#�X�H���ǂ*��)s׵��d��''���$ }�� �S띛�21Jg����1���:!m8������U���8g���|W
��n��F����p�&���O]��1%l�s�ɫ�@��(z�
q��Y�*�*&**<[�swm�C`)�g��e�j/�8��#�'�c����<΅�o���Ҩ���x���$����7�bl�S�T����J�'b�G��o{��`��8�i�=�3�`�0����r��9�Z�ѧ2Y]�>�h� Ia�K��?7�w���F	��K1������#V�k��7g�g�_�K�|�ł��m!���$J!�l�v?ФOqv8!׎q�����ws���ef��9��{4*,�*6ob"����]�p�$�JY��(s�K�^�?m<"/���@Wz?p�lm�r�����a+��]��i��.1
׮;�X��Va�:!g�k*�ŵeb�0tL�݂��A�'(� �s�%x<\%vX.���Cy~�9Mp�8��EU�m�]�m�T�c��>�!B]��T*L�e����1���᫷R�g%���ut�����_���a%��P|F�"* )L���щyq���v�6�u%P��"6w���|'�5$�̛�RG���Y��x��V�$����A(�z�Ρxs�^�V�3;�+G6�J��B�����-\���5����AX_���j��*��9�S�?#�UQ�L��HLa������y��q &f��tsZSW��j�l?��?k��R�~��'�zJ�3!M��+͞aѹ����pG�D{<|��M������ g���;�}Ca�8��s�����!S�O�қ�@>{�������g�J�pX��B��vƭEL�>�����?�CJ<���X�uK���f5����;���e�q8|���FH��QB*>�q�f��,\t�*J��]"�Z�#ֲ�qI����d���&y⭍�Ҁ�����d����kaM����I�6�u%x�+�������*?C�/���?:W��d��Ko˲_p�ݵ�rr��-(�� �<:�6b�ua�W�m�`?��"5J��˾����Gy���D�'[��B��}7�/1CF�Ph5}�l�R�d�H"��L5����(�) ���GTl[�
���;�-!}�_���,��FJ��OZ�����QA���)����]�Q�Pv%�F��#Jg�UYm0���jӗ%Tm�ȷ����i������|����Kn�3���̀��b��&+#4M��+�L����1Jw�h�Q��	����{;���Uܞ- ^X�9���HLr�;�|V�+�R�j�ب]����M�/ij|+d�#u��J�={�$zf�6o]���o$禎��B�(�2�����S��n��,�{�s�L;Ao�!���#���P[��d&�B��VJ����Re���9�i�tQg��߃�c#��X_ŴLOU�ϓ�/s���n"=/h ����B�+G�Ӷf��x���T�u�l���!�i�#�﷯�v������BƂ#Ԭ�%C��(���˯���$��h{O���@1-�zc�Rwc���&G�R�Q*����1�&4�����>����y�Y��xt�U�N@7�d��̧�)[���+���lj�Q�lo�nv�ο3}5�$�*xsU��.� 43��=mI?2�?���oD����c�j?�s�2b�]�ʚ�*�ӓ�d�w��:B���gw������v��["�: _d���I#��^��t�:����ʁ?�cޖ=�3�L���<��3`��]L3%D����-:�U��HS��Ê�R��0�}r��?��Hw0()x�(n`'���
*�D}�Йmy4��bxO������w��R��̑:0���wL�Wd�O���� ��h �ҋ�j�w{gpH�ZE�������L>�	��@C���Ӆ�0���`{e�e����|�E�{"I�V|8���5��Ϸe*��8��q/%���du�@����!��O�_���B7*q�@T���(Y�R�W^��ߝ|��
�1،NCO��~����@ۖ!u��$h	*����}��W�N��eA�"u��C�])/-��ck&�Y�M������*�l��H��e<]*O�i3�"&
����d7۝ݿ�NO�u.�GA8h��#�����O��g��Y�}{4o]�%Jx�x����>���.^��H�OY�g�2�� ���|=m���QO[ܵ&�?3g=��f�o[|�<��'��{i]���X�vA-nQ[J[���ۉ?�#����/?��	N�����
��U"�Y���Sq�h�~��Ъ�ZwZi�N$��0�v��@�&�Txj�W��v���֬����$�Yv��^IFs&p���N��/ ^(�/�D��L٦�ȩ�Ç�IH�_����XHM�Հ�:w"?i*�/���1�m0�wl���;�T9�P�>#J{Wҵ�����������C�~~GQڰ���?_eK��$4F;\6�Jf�5t�nܝ�s�j5؞;�eO�f�Y���\�R�V�9��ג�� �Fj��,�=�$o����$�Ŀ��T�V6	-ir�Z��wN_��'<
;��A"�(c�޺��K t{��T\׏p3F��:#O�7��C`$ܐ5�ޏw�FKo�l��9tQ}����T�s��ͭ��%M�.�UѪ}~��{�͋��Bj��V�;l�� )��#]陴ck�q�)�f:9𭮚��Ղ���I����ֵ�ĂR�$����.�t��of��Ji���ωH���7�a����qx�O�1+abYYihbR�����
ed��)[�����ཞ�]ki���O��b�wk<yx��L�lEN]Q�8��}���:�tf}�nĄ�u����u���X�[�<sJ7`�\�Cݥ����ÏH���[q���,Od��_�o�_�`�סD�]�1p*�qh��l�*_���W���c�PbM</iFͩh���˵�(2H��043
9~�v5=�l��yr����U�����s������X]��-٬�W�jRC��h�%�K�����I�ݮIl�IT�O����ៅ�܄�����AZ'��ܕ+~����M�Ds"&�~%�*hO�}|U�9̈����������p'I��@AUxo)S��>m&����6�wz&c�%td����pGX��5�ڄ�/tn�v����ٕ��OV�0����L�n�ϐ��ک�Uh��HN��M]���
a���{@�7�%R��Z���;��ܟ���q]�v�B�j�f�r2�a9yݩM.��O���c	���W�&�VF�V�\,b�2��9K̐5���ǖ&�I&4���e�@���&h	��U���`��6���T�&ells�(٢?������3�����'#��}#啀%A4�nGW�**���Z2T���_�2���}���p�w��F#)��� ���2^���sߕ��u�����[���}��t*���n׫G4��I���s��s��f���@�1�sQ�:�.����GG ����lg��Ǻ���&O���a���d��ֺgY�7pf[o�E����TDV��K��m3�Qߝ�	99��^�伬>ώ�d�<)9]�������ǂee�x�J�n������vvG>��	���H!'1N��i����)6VZ �h�9OCs��!͸ g�L�Rϙ��ګerH@��	�i��!��J�����2��DI��A!��kŎ>�C��'
�wT��HI�j������:
�`�'�Y��A΁�! ��O�D?Ta�Cb�U�/��u�P-X?��imL�j���b���| �}���&+���{�Z�ܹ�@�,hE�"�h�p(("�����74��O�#�\�u#�����
p�1�X�&�B?� Uw�Ɨ1o�`���4�z��H�����s������z�*0x��<��k����������}�~7����{���l˾��M$������9㷨�Ó����y���/iB���b���)Ao4��p�}�ݬ���o�]�~ip���	��)�1Ld�C�No���ԈW9-#+h3�o��f���}��g+|���xڸI��]}s�t��tt����������=4���;�o�l�E6A8��Ж.ގn��h!��/�W�@ A��E����}������Ѐ�I��L"�T�3/v`�yKڳ2�I�ILca�����q��~�􀪊S�MOg��Q�]AR��?C}���<�!rCy���7�Rtq��/lu��!�G/�yto]�����n3�ă$�)�����>�Q��j	�iu�� �
GGjP{[a�)0F�򧼕I�hsMsn޲�����O���pppBz�L�"X��)����x#����WAN�:V������A*���N1����z���|'����]�����Ӵ���T��U��Q�jtb<B�۔S�p{�����n�'h�_!�=��,����pX���-�o��Vs��x���~��ܺ5� >�]�W$�Y����M�5�dZ�$�ݛ��ѱ �S̒������)㧝Y;�J �vW��Ho������c�Z�&���_��'f�Tz�Y��T��-h�����d����~����:��	Ӌ�� �͇X�r�-	!%a�+w	���k�w̴�N�*����Wnb' gL���T��Π�j�֛I�:�|0R8����6����Me�=2�?���D���o�P��,��jIm���T�����9���*թ�:�	k�����x�$zj2�S����pgf�l�s�Eqg�-I݌G�{O����[�HL�L�����y�����֫��ￓm��;�L�A��%ER�(G�h����ae^��|��T4��u��b��^�;������ਪ�WT]��\��M��m�[�W���*_!AyN�黌�τ�(�G���oh���>yOt%�;��\44��3�BY��������º�I�=��x�nz{�Aj����50���5W�A��6H����ů@��/��u�yO����12Qr>���{v��<M��m�p��=��������v�nP�'D��4�;�Y@�D,"zG�]�Q��
������/&4N�)�ށ�tl��=[���+-�[�o���Y�F���`�{߉�U��|nN9k�B�)s<OE��u[��cP�l�\�Mu����y���x�w�X�<ަ_��YP&�+o�<��f3�,�0�ӳ|60��m��(R�bFm�gD+����o��6/.��jzi-x����glі�`��3��:�/M%���?za��w_ӿ���ˊ�Ꮶ�~ɅQ)�����������L��[{U���{������s�������gMS'X�UŹs����J�1p1�>���V������cvZ����C� �?u�$�-��D"64���c�ZSj�U����or�(��9��Ľ(��f�`�����]'�n�����:�������C�w`���A�f���&�pZ���cE7��:���ۛ���9�`��$ ����fUڢ�JJ�~���Z����ۅ��}9E�̶�w?�q?+��VT�jh̫|�oRЂ�6)L]=�S�N����q���:1�':�pM��x��@sC�Yu�#ŏ���.�Ԝ|n���eE��A�T'qF��3�^s���� 2���o���	s�x>	����ע�E�fA�5J"mlg���vn���s����kr�@�er�֙�[����[n��^�	���;�u�|X�[�"����	;�Y�~�8�Ul �����9RzqcqQ3-�τ�Xs�-����%t�� 8{��4�h��pիS���:*=p�.&��)xmzr��9�����d�:߬��@d�/�5J��T���t�Q��l��fw`y�'���R$!ŷ@���g+��S�g�a�5!��FU�2����a���!F"�{h��ک��/Ļ"�{$Kw��qM.$��'�u����ٞW�X��W���5�Tu<��@]9��x�q$ѣP�d5<J%-E�/���ܛs���4$`�|���p�O���@5],n�mBI����G�o�q�l��Y�� ����Bt�/5��3ԅ�^\��^��J
s=R�:�Xڴ�?��d���]F� �z���H�h�>j��?�V�Gb=m>�ã���<ca})h|��֚�
;�-r�3~��1�8���65�w��C[Ԉ��#�}���5���Wf����E�P����ܼ��������"SC�L�����^�MSl���7U���ízS�L߉E!q���u<��I��?șK{B޾#_�b�O|>q6q��a�ckh@�s���-/� m��˩lU=���#�����m�%-�8}�2$���yr��}�4,]��s����-��lI�y&�}S�<5�����
�b�r}�R3l.��P�m3C�*a�U6�&�:�8��58����i� �Ȥ�H󉨠;|�-w�|S����]�w4�1	C �Q�џ6�ur��HJq�!;=��lン�u��$��<�di��}z�b���4��E�y�P��nψ�����	��R˛�,9^a�W���{ZA���?�V�.��N�T�?J�,8X�fJ�R�@t	J���|}	�I/��k�??[V^�v�nd���l�Y��5��;���̎��C���ze��&R;@*9���ͯ�kۆ-Agk�n�f�����Ŕp��`�� 1 ��Xu�t�4�h���U6�7t�Slh�#�w�-M�9����Kc�T.�{������G�V�[���ﱎj���w�c3�|��������+������~�>8�Y�!�FC%��m����q�;4�&��� 6c[kk�sc���|��U����q�_m��hlۏ����c�|Rٸ}c����l��#���|�moS��ԝ#�pn�H�!KNBc��@s�I�VvV��Vm[���7�x͟ ckz�ɢ��r���
�TO��{}S��xmxY������f�'��>��v}����A_��x�_#��9������zԩB�9l�ck�^����NQ>/�9��F��WA��7qF�����S��K�d��=���*G6=��!Xݕ���]?{���]k)�ͻ�ƨ��*��̫d�p]aX��/�_t�E����w�!�����gf`[�(�ҩ���zČ�4��@=^u����{�(^��@�~M�Sa���c�*���r�T��z�����-�FCx�˳MM9��������_�i��r(�A�\U����G�<jZ���yd��n�!I��֖���G^ytJJ���i��9���ű'Y-�$�~�����EF�7�֘���vD�M���I��/������~�j3e72���Ë�5���OZW���Z��w�ۃ�^�N���v�ǔQ/TA�x����=S}��51:Kp>m�>ǏNtj���_sz5S�<�IQ,Z��y�m��V҅�+������?��iQ�m^q�&x��m���Ûda뤾b�&������7�2�&�����̤1�� n��OhR���T,������04>�I5IY���#R��D����T���?2O�����\G�����H[l$�}L�[�FOٜ�B�6�i^��������䓓���=x��ꞛ����Z����un9cw�Tk+��׳��ϧ�P����������v|)��1��a�-%s��y/�5xB��(0#�e�B�Ɵ%���=E�ŝ�����Α}G�
5l��	�����G�J�x���u���/Nm������GMM�uDkY�w��q�Etu#;����Z���׽���D�I��u܋V7}���5v�m1��&y!8cJ��w�-��,�8����O�f����;y�]��=�7��E�麗aE���:^��%U4.a�eR���Y2Z;LC�v�tMeq�$��I�D��(�bw,�CJ�ö���r=`t�#�g�(��$Y���׉��d�)+h`}��\�.���ͼ��+�:n��F{9�8�0�ؖ�n�[�$�wUtm����1x/�}%��s5ۮˁ� <o�q{�Z+gb@Ѝ�\�U6����=���w���� �@9S�p��;Z�-c��!"��vᜁ>��'%���hp)��p�o0�`aW���ho�v����.���-x>Ԫ���i���}�.�U3w*|Ը�
5�c~��V$X9^Mp�3�j�E��>����֍�;��<{�N�#��kķ���F:;��iL�I��.t���G��槪��*,踬q��#]���ย�Qo�h�9�S����CnV�!<�}_�.*>�����} �w��K��E�7���`y�f������bRedR��쯝�1g��y���$��(�
!ͮ�O,�!R?�@��/L�<�j�n[���@Qŝ��)L�w&��wz}��oC[cƗJs��~^�`55No�͚z�7��/���1��e���7���-��Cu����(�d�~��r��T�!��߱jJ(����M$��]�j������F�ˑr��0+-����⤣�~&�2�������$Y��ۥ���4��P����8�����'�g#��{=�3�E������9�^i�`����������@7N��(��|��$>OVgp9#<T�xgzk�K�}��M==�U��)̷���3Q�Bk�똌Wt���_2�b��.��	=�3)�^m`ң;����j�4rS�K]��\��M�'�����7�/d(��& &{�-P��]���e�k��RJ]]��W��7#e��� ��vt,ʽ��x�E�����Ҭ�zV�C�^[	�5.��:hqN8k�`̽���O�
]{���@\9�Y�����C��;R�ORR>��/���z�+���70X0�m���jb�+3SO?�~�v�ˏ;>!�I������{Oڬ�[г_�3A�X$�L��f�{h�~����1��r��c��*�'�Tg/bk{�� >�}�$c��«,	�X��K����R���nP~���B���@�el�!�e'Afb����۷���.e�D�ï�P�2��)����P5��O�)�tVbE��d~�Q�(�e��kNp���? ��
��η�˛Z'w'�y��;3<��}��1��Z�:��|V7�x����&z1�C�$����C^���zI�qN[AmW���a?��t'2������ ��8&�}3�*�����?��">��宑]C���c���)j��lw.��䛛��g{{k��Ƕ�����y��=�`����쟭]+��)I2�����cMu#��	[��`���<��[5��]E�y�R��IH]pڮm����O-U��G9X��o�sPB�e[ŏ;e�5�@��
��?6���\�l4W�:� >�%\���-u4�#f=_�Dr̽�~8WB�N���8��?�hߵ�n'�%��(K�ҟ�GBv��������E�{�|�C��3g��-�6�k������t7ǋ��zcO�r�۵-3#%�rd�ئ}>JArD��J@^"���mj�@LibLm�m�U�,�
?H���������yb��f�����zr���ߡa�ٽ�n��E[��T $�����Y�ȥ���&���.��GV���W������@�~���U��
*���f�g�+��@���J��C���P����4eJ}�S��̵��d����H�FGt8��a!������3u$׸e���/&���b�c�����/E����*?1cd]��� ^�^�M�Ÿ��A��Z&��J�9��#�_���~�$�Tt�	dP�v̠]��_���g�SF���b������!�3���e����ԸO���ۄ��-�f��kP�ӷ4�������Z�9�M��T,n>����btB�v�~%�{�j���O�z  ��
A^���7�{p���UV��%��V ��w�iS,
qd���aP����s���\����M���!E��JՇ���O�F���������#�d6�sm9����r�l��&%�H��=27\$�cf��v�Be�}@�7""�2e�/D�>���Cv�>ܫ��cMe,@�5���g_�0�s����5���=�AZ�Aًx���-n�]�v��'�Ɠ�`���-Z��dB�N�����/[I�'ۄ�`/�l��Cb�g
��E�c�Vt)��mǦ�FK{������3�?nވ���{����(����R\̈́�퇋D|�K-�f��#G2����]�	�x#q;Ƚ77�Z������Η��c�?g�p�/8t�P��U�gg��[X��!��ZY�0,��;���_*Y7�|{�"Ԩ����FO̅Qr���5�l�+������2o�*pSxŖvcx�ه5�G�ݔ��W�:>u�䤕�$�����'�����iB�z]��s:xƬ~�_d��"ۢ
 ".�е.J�onib���Ж�_�i�S�����[���7-M����pȔQ���k��|�J�/�j�M�
/|�9(�m�[b5^��s�i�Rٹ2C�C�+��=���th���d�0�$1��L{����lYĺ׿���T3��7�V��˞hTʽ�0c��]��������5?͒�ˉ��%����,�d*��N�hy+�q��j=����>���Zc��1f�O�𼤩�0u��R�_�أV�{t$�gTXGN�ԌW|���Z�0�U��q:埊ff8�Wַ��P��M�4�UT[m�6�w(nm��P�)Nqw��;w�E���C������y���'�$ɚ�r���H+K7���ZI�b��2����\m��Q�2K�<�Eͻ������[q�uv"W(6�\�?�{c���Vb}b�!���XY��M:79�(fT���?*��Tä����K���Z6�5��ڋM�s��4r6Ǥ��{ڵpB&S&
hP����-G_�%=t�(5"�@Rõ��%3��+�5��Gk�n�k�\[��N�Z@�f�T��	�F Ϗ�ݮ���=p�kFR��ϿXw�`R��q�)�zS>��K2���Tf�����lY�����CG�*�O,�B'�Z>�5	 �G[��9_��}^pà{��EH���ɰ�t�Wwe�K����	b��$zY��E��R��{n�#�KǞ�ڋ�s�>�%�U0��l�f�x@A��K��S�xl����� |5��֣ق����ZG�B������z���:�F�5��w�N����K�nv���HjU����6{H���Y�*�'7�0#��u��G�Q��e��.���9�1�NWg�!�����4�`��,[%���Ǘ8��oڦi�~U0e/4�U���vj}2	x$}�~ژ������O� s�Qe����
N"��������������t�r�W~hm��I�b6p0�;ƫ�p���������_dA����='lZ�^c�%5��p��w�Z1#"����ůD�!��1���j���Va�Y���Z�B��n��Q\@B&M6}��խ�8š��."b��_(�e�Q8��+��K�~iw��V�O�[�ZƬ����q��5�p�n���R�
�~p������5JM`�U�������2��/��R=�]՗��j��b@��F��3��]#�D%cG$��f��	�7WT'TV�]�zE.v��C����t��I��A��OrkY�&X�V��nV%?�¯	���S��⌴��0��T�����3c�T��4�s�k�9|��ʝw��~f%c�ra���X�Qf�\��@oG�p�Pj��!n�8>~�acZY]! ��0�~��v����,{>�|.����q9Б���ﲴף�F�m ���w*>�p�B�W�[���v��h����*g���+|�J�z>5��q�-�\o��}H\T�ys�
�]��m[G&�����d��������@8�޲�&I�X��� :лI����3�N��d"�Oh��+�.za*��>����|u3�B���zCW�XW�Q��[��Y��߻.���D�	Y҄�����W�����m!�W0D4ȵz�AZ0�YR�>�]�>[��&�������(�*]x�����%��ܪP�@�h���T��������S�K[U��'��ת�/��J}���S���C]�>	/3|B�ԓ�W�r<��$��7̯<cQҤ��|C^yK�)E�eR{�� ɡ�U/�G>.�����9��O�������$|)jcs>k��6�ADE��8EG�	`���}d�ޣ��������6H]{bl�����Q�b��к�)�:�!���^�A�3-�5�n��s<��q�v�g�ƫ{n�y�����ik����׏J�	��]y�%k]Xv�b���U��q!�"�ߙYI�}�0,��7���w�x�7��I�)E�PlTC}��]�^�2�����R�iU���G�����lD�fE+�݄�0+�,��bW}�\ %�ã@�T��.�Mݿ,3�)��4Q��	�.谺+15q�be^���D��t{�2��6<���y��h ���mm�:�1mBظ���O4�f/�),�����D#C��] �х�������"�rAI���2d�W�
��$*(x�;5�"�	8)£g��>�s��3��t�Q�M>�_w���rD��q&4�c�����o�i�77�h�fόdjn��!��79��,���uq�|�>+��w�^z:~��.���܎�!㯆 ����q/"�k~3\���t2���#	'�17�<V������_}��a�!eu��@ �ؿ����\���Ɛ�3*��_�����ښ���o��*�{��&x���o�iP���:�<�u�������sT���`n�����9n�/�.��50���2�Q9�]�� �K�|mc]a?����ug�o��U�w�1<�Y�W�����b�N�qqn��'o��j����+���ũ8i-�eGzH�ǲ=�ݕxU���y��k����'�	� �r��Z���G��"|OM��=۵�ҝ�f~��	:_���]U�K��~��ɸ�ӂ<8\�-fa"�����t��<�(�wRN��@��HV�v�\s��\]�Ɛ��_�:�Zg4�z;�)Ύ>�M��V�� �y�P7�aX���2�)�=n�x\ƪ�Y=.�-��	-Cs��}��%�J�����"|n���C5͙ɿ��[��p�U�L�����N�ZT됧g�����m��f���T�f۫�R"�y��/.ӑp�~}���_�g��l7�3S��� -'R�ۗz������'���#���?�ZuwMDo����*��\�G��JN���iޅy�?����ä���ҥ
Q�O�V�E}?�Ed��w�A��+� ����:�1�$Gp��&�l��BF~�# 9��@,5;���#[[:z2P4��b+J�0c��	����W�~��5����s�&E$�� ��?o��^�I|���p0�
���G)]�@]���j��w�&�߻���L{3݁���fo.���Jzz��)T�߼�Z���������1Κ�G��RA�q��0']g�P���ڀ�+ߨ��oe��	#C��J+��7@?1ڳC)�P�4�ؕ�	����]�%Eϒ��&t��5y��kf�����m�q��mZ*���!�&v��<���8Ubgl�!�"ν��}~�4�>k�ՃҴ`�e��ƾ_���-��@����n�Jԝi���6�� ��Cm��68�!�£ֆ��`�=n`�$U�*�����u��=��Z����y���Kh�Z��[��¶�yT���$
��d&���	�~�}�D�'�yX1i�ֆ$*���|X���ي�3�ԏ(lz�M��wǏ� B��+ڀ�D-�v�!j����u�^����<d2�����y���H*�u�ƫv��B$�����\����U�IN:�QX�Q]<F��1�G�P/�'�O�>�.���$%\tz־�i��^���7*ZD�9����q	;Y��y��琍,�F��J���w�wp)��D��O\BM��0-�Gx�o����C�����z�9I\:uZ��W�߈�َ�y�X%�>t�����u�p���X�6b����N>�z��*��eJ�|����N��ۋ��
=O�����4Tά�J��d v'�<��E�ZOb�K�5]]e���%�	��.�]q�(���҆|�L�9���,�u4�BJX�T���)��&@�(��7��AW�<=�/��"DVVm*��ZbG|M5z��-۩ԋ;�K�]�x>�uy��Jغ�}}��3���&O�v-� ���šY�g�?2�������I��&c�TrJ�J�����'�,e,��e�'�곝P�j'˕�s�t?������	Q����5[�;��%��\��Sf���Ӗ��N�H�18��A��I��<=ظMps[��yr�J.NĖ�:0�c��LS�v6��a���0~ ׻�����^�	�H���rg�$�ƅߗh%Sb�eT�&@�̳sN|<��*�ꔏ/�Ϊ�	�ӑaQGeJ4�j;���:V��d��9!��b�SIAl�Bs��dj�_��*�:��l}v�hG��4����k�s�ݨ�%��S����LȽ�HCo,d�i�@}�:�}V[��-[~�h�;cv�:�dB� �gKEo�)�l����#�����+aÖOn�����P�(;�E�W_�#.F.��]��|c���υ��P��� ���13pl��{��1k&7I�=�WG����BN�K�ʧ�j�كwΝ?�+{%P,�j*/��[��L��8�N��������>nR�6���e��I
��y��~��Huu8be����L�#��۪��)o����U`���6�z��qU��Z���.Q3v�;�6��7G쫵h����{�Ŋ�E�L�}gS+0]5�A�n��MQ�K���HG,}��/�x�zY�jh*�_�27���~�(Kl��#�{�(Y�E�q�WX�e���4��ND�5Mk-�]�P�g��\ �Y�Kh����#�侧bP��+\N�`����7R�V
���p������a���mYuC�9��"�r3��S��鎋�(̱I:����D
�!'�B��s�o���A}�׷{�JD�ޛ�/8�;�u���Ĭ�/}ʗ�3.Q�n�q4�`���h��q���r�\tҐ��u�O�úgE���@�E����kM��m�2G���S�'��_���l��[gi��D5SĨ��QqD�"�n�'���+ �u(����D�0$��"�<��5��vr'�twL<g�DK��px����HK�7��eDa���/�8g�m��cě�gβf{R�=c,�=��� �ʶ���o��r��?Ɨ��fE���&�n���ή�|���46���SRR�ijr��'M����E�tja���¤��X+,�����P���Վ��]#AI���b�����]ٻ��_�o�I���4fs�U�R��ș���e͉/
;C=�2�$.+�w9��'^�����V���d�!]��ޞA@ E�����`(a��.0�D���OEO0|۲��:��݀[�Ӳ�|�p�5Y�E�YZM�ܞP�]�p�8(2�4m�[����֖5Jd��k`����D��-��?5��6���Н`�s�;��9�b:�(|ս�R��]>,/�z����Ý0o�wu̓�u8�GA���I)��[�y��
& LZ�!r�c������}I���B#�>�e&%��m��r�i����/�H��N�gaa��9��?������O��?���{�*����@�.7J8�ᘝ�8�KK ���9�(z���� ㈜A����3��b|�tQYC��D7Z�&&(�)�ěU�������0,U����bx��N�$(�t?m��iO����	�+�	���U����ɌDm��>��}����H��a0j�"BX��iOX��0ِsp��h��G޳>������޿5V&���~ܷۨ�g�n̽\.BUh?�wB<� o����ܐ�1���+�r˜	8kݱ�FLNNwp`�W�x�q�����Һ��1ٕ���|�k�^����\�--�p��p�IIl�DJ�r�����Fr�\
)n-M��U��| D㾟F����aY��Jе��a�+j�>���_Cw@����?++r������o�N��`��$����qcjxW����9XB~:���ggˈ��КI�re��?.���c%�+�s�<�|��Q�{ꦦ�տ@	x�&6���k�}(sd�^��mow����5�r������ ������Q�ݐ�x������W��0?뫖#eT���WG d(��ҝ��zbO��� b��}~�##�)|����Vh��v������콧V���o�������Y )���	�=~�o[=-��C�(�)Le��e�6��+u��[��������׾Wk��ҨN��À��T���һ��<�EO){U�xy���L��j�r���r���Q �s��pE��t�/�2���]����\��빂I�Aƃ7�`c>�_`Ȯ�t70o�C�A������;�U���=�}|��*UL��ֶQ��l�b��0�ൗ����r�׽F�?�,��?i���@����m`r�(ߖ�4�@P�R�B��?+�v���7̛���7:�5��+��v��n�򻮢3��yUI�;
����+]B+���-p�,��7�o�7��C+j�9S��d� �#��_����s�S�1mn����Υ\��z���.v\��Q�!�����;Z!��W�^$K�kQ�����0?�54��1c��� sd���9��7d��d��L !�]�O�!�$�A���_��N<^҂(��Bi�X���^�ߍe^�Bj���M��CZ�L���0�(����;MD�4FءϕɗV�L�ð����~�F��bZ-(���4�`��|�.0��e�Z��9u�C�Q�2�GC�L&�{��/�y�IH�,[~���]�ǕȵR�'�1L:L����ð|L˺�H�Vtӌ(�)Vi5>�Ln�t@�D�!�r�tM|����½[�����I���e����'��{QK.�pH+����=��^�%u�|�0:£���i9�U��]m�D�SU��q�)�%�
��|J�.-sYX�Me+]��TgBN,�_������0�C	�B��Y2���������Ta "�3r4`~�#�O`�yұ�.��񴼍��_�c*$�<��&)��)��e O}|�͖CZv��(oTʐ�j����3�WKL۷��|tc5M�2��Nn&����T>�k��N���y����I��T��\p��m$���I�nn'����!�FS�nk�=1�;�2������gb"��#���~m�rm�P�gO��Oǥ�YF�[	�:}�/���oxӆF5���(.�cY�Y\�O�������Q�\ou	���Y��
 ��]��{>�)IT2�7e�]���VjY�2wW�7�vv� o�SWs�A�
iv���`��
�)��KF�i]�e��a�D'�pmR�ۡi.�:d��MhoK��@��/�gj�V)')v���yu����hPNL(1��ч���tǙp;�>tx���qu?x�R�;Kq�hyq{P�1Mef�f����7o?�k$Y�����W�BD"g� d�����1�ߥQa��_�\�
��\d=V��� *Os�<�9�SJ~hʸs%�/մGV,�o�ݐ6��?�|N���+eM�".���(�� ��둪GtL&#�)����<O� �^Щn���07�K���CW<�R�@9�v�s&6X^�~ ��ߒ��f���4D�/ �Rr�)ڍ�ܘ��y\�4��Z��M0)Ήв-H��anO|�ZA�;�l�W���Zv}_�W��ˎa��D�_W��D�*�XM�����I����p<���f�&��o�kqm�g��������STX	,�н��zL#�3O�__)��f&���U_���n����m\�W�3��gC�O�0�J���~�5G����ꄸHF�mV��/
�|�6�KҨ)~���	�����!M����4�@�ﻛU?��OB�'m̕�8��������O�\�q}|P���H�S)�O�	1�XYR鳆�$�K:��nr�7�P`QV\�Y����^k�1`���ZgN��15c�oӸ�U~�r�U�&�m���t��!Qb7�O�|�ֺ�\�����yOj�;�p�buu�V땫��-��#.K[ڿ�Oj&�!��� �"���qAbw{�-��c����6��,:Ual���dW�]�8�s�㸇�<��L}A1��Fն��pgn�	li��?0�50xs��#�����Vf���������ʞ��E�.p[�j<2�&�oo?��{�7,�@1aX��&aA����su�Q.�׬E�>l��x��-7}x�vޫ,Z�8v#lD�e�H4��u�Ne%{��g J�*�F2�d�q��'�^Q��L6U/�=����M����$�3֟���� �]z��|��\לT�JzD����Ϣ�\���R�Z_����hZ~��[��IЌ����7�bW����/z�I�K|5�����'6IDG�(kB�;�>��!��7��
�����NK��Gs��l��&�_��w馑��/m�I�U�Tڀ�t<n��'��p_=������x�Qw�.9};�EC_:��uX�w�z�ˡ���67żn�i��m���E�>�x����ເ���>�·��J��e+H���N��V[9�g�R�a�!&����	�����ڣf �qb{��=� �:'%lM��	$c1�Z#����h_~�%s�п�8��~WpK�I�P�^i&��x�o�͉�O ���}r�|Q.F@i�3\C�AI��_��@�a@���~P��n>�k��lԭ��`G��]��5�N\�qM�k2��ͨ�3�������CF�����
�Fo�䓙^��L=ۄZ*O^M�\�Et`��S��W����'��GE����̓+����Y��M���qzHas@_ao.|��AB���>��	vT���+w೫��;�����w�h��U�q�1peH�2��q.u�}��Y�(���c��(���4C�z�B����q
��������K���8L^>�NS�]�e�j�$|��5���Ii�Q%��@n�M�������M���V@�Ii�X�5I�z�g)��H�R�J���ڬ�e���r�@ҏ�s�r�kM-��C)a���Z���̣�Vkw�+@�|�@�փ�ǲ�H��J�U!��9�T��e�,���B��HX��	��k1_�$G:�5лu�d.��O��8*J�P�˗��~ڛ�s�Z�Wk��곇{z�W� �*�+��Ѝ��X�c���w���}�4'S�G?���Z�I�U���[��}��e����zJ���}P�ě�2q�S�d~ڛ`œ��I�^�4���ZH��>`�[���X���а�������F��J�$5��� �c��>CRa�+���������V.�6n�0�Z\Ͱٻ�w7��}�ɦ� �8�f�3��ƾ�3[oO��@g�����X�SGM ���M�V�xh�xڟ2Xi��h�I���+YJ%BvMu�X������U�lgB�ƫ�ʤoB��
p��<a[;~�O���D\u��䄉�=���n��xx�֌�CG�l]Zfw�wF�k���+�~��4��e�����Xi6�J�+��"ċ����fo��e.�R�chI$�{j�����;+���I�̳;q�%���5���n$	I�@�z}�NH�^���:�`��7>��=�83����΅��un��~ :=�a��!��E,�{�el��ħK������W7! 2�T���>|&�h:g��^o��Wk��Ã)�%�Q�|4aX��KH� �h�)�Y���%;�l��^��e`�i�!�#It҈���:�׾�Ͽ7�Z6댘||��E@Oz�3{o�5ˁ��T����������S(��h5�!G�jͼ�Pq!��1yo~��H��*<8I|�����������EG7l�2����/�Hda����*��/��+���	�FX��8ɷ��� �Ҡ^_k'�U�iba� H�]��	m��!��`o�=�<u�R���=^�ʫ�e������|�Q�%P��lwsĞ=�D�Ef����]�fB�g![d�g1���h'?vI)-���ӻ��iK�?���W������<oo�$�����L�O����oZ"wk���岲!F����ew٧�ӫ.%g�&�BG���	�������k=��Z%ѥo��Aů�C���㉬����� �5SQ+2tJ�co��Y�̣ZG�����3��k�����]�i�T ��*���������>�$�B�p/���,p~�h�l�_;|Y�J�w���(4g6�f ��X�F����yr𞒵���k>ך��
k�kG��S�<����Rcj��]�����}�)��}f�ʽ]�I��ϑ�Z��W��8(��}UfX0�&O�=�@�vAN�/>�zϽz]��U��%�U��TKd���y�jQ�\�.m1�����]�V�hot�V�@���Q&H������m�vƪ뀟ҳ��yx�x$o�7R��w{ۻ!�ɉl�O�����{��7aeF�ٮ+� �G��_m5F�GH(�"��n˸�U�^��'�껤"�|�{<�Ar&(i!m��ـ��N���Ͽ2�T�/�"�.��R�<L.?�_HL����<G�p0��QK^��
�Ǆ�M߮� ڂ ���>G\��?��*��U�}�6�or�{'C~`?3��rt��s��yο���=Ii�����a�j�v@0�� �Z�s2�WX��Pr���HG�4�Y��t�Jp�H�<�.K{*P+SNۊe�nEk�q% /��7��c�c=ݱ����۹z&�����@���r�;gl-� z%#{ �x��h3'o���#��iRrĘ�k�$�Ut�n����.��E��TPa	2_���K?��L�|�?��WI��RZ�r��Ɩ���	st|sU���+�����I "#OKG�b�X�lC]�/�t�%�.��(ԗ��t$/w�s�ѓl�޺�}|�x��v��ƃ��,�(YU�͈O|
 �e�y_�xΛϬ)�o��᤯��,�ZEn7S=Fjθ�hf�_v�V�=�rT�����O�sn:I�H�i���UT@���>�>߂�)���Il�@PDj���.Gcvl"K��m�*E|�WEM��t(�����@gR������wa��N�ߩ�O����'vv����#~.�GaC�yi�cr>_�}��A�+��MX`\f�$�ZB�▌j���"���i�L�4���D!m'M�}��C��R9�G��|��Z)"v��?Zm�-|WR��S����]:E3
ߝx{"l]��!�,n<���RJ�0�N�U�&�׋�,�`T����h���2��S6�d�o���yY����5@W�*\�j��_$6�|�w%)Xl��Z�h��Q�Y'�ϭP:`�_q��H�fGz������̬H�+`�����kp����f����񇳌$��p ��m/�|�e�z��Ю���F�.�G�H>�g9����3!�1T��C�׋�U3���qU��_+�ZeJ9�D	!�itΜ5���J�����KOұl}��01aId�in-ƼKT��d�M�I�����cֹ,{���]-0�c�G�R9����*b��ϣ��&�~���":�7M=�]��I��Z�5<|vI�|�ymUA��'X�I��v0z -�mĖ�V�˻�mu��I�����=#�:���)�'��$���Eika��������f�Y>��פ���Ë@٤���I~]2� �Z���,��?s�'C�|S>�K����`p��nayk�ё���W�����X��b�6�x���;���O��KV�Ubͽ�e}�~�u�����Ge�H�)��Y��up�c2"��:�3W���%��ߛ3h3��ڕ
�i~�?^����L-�?JV� ��s�)�=�&0�Bu&B�õ�P��k�7��Q68p#�L�u���#��CT<?[�:\�_`lA����{s�9��p� ���K��l��U���%+ӗ_��{mlюy�w��Bv��k��n�m8g/�]"_/�'��=^��'u�2��5��u�$B�~La���u>�k�ύs���ŉ�P��{��^G��ƚ��3�|�b�_v*�`�Y;�u~�n���~�d��T���P���k����xs�E�
&�n�o�8c�����_(�x�cv�g�˯��d`��C��S�kz���L"K��������/n2����"m���_���:;7$�)
����BQ��0,aΰ��0w�ɍ��8�v�%�}�:7���~�}er�h��t^,�8�"��/��7��{å��"��)�&N�敯�ןw?ù�k-�? �i�Qu����yj%�?��D��u�њM�ll����&>f�2��z���������|�Ɍ�bx�ƼF�Y���R1h��I�]�Z.w;DN����6�+Ƀuv�Bd���&rӇ*�ɳ���xƹػ:��sG��Bn?0�oB\�Ͳ�nki%p�V���Gx<8�[Q�]f?1�m�R��$|��>�<k�p�[+sR���	�\�[���}���_��R7� )���a_�b�|M�g���(.�KPd�O�K�+�%��c�|[W��ɸ��ˈ�rR�B&"���\<;�Sc�������W�8�O�F���N�(R�[1����;�d�SL����L)�iPo{�V.���](�X?5�'%^�}�ݿ��NZ���>*�T�Sy����}s�����+���Bz�H��mkv��?���<6�Me�|��|����`�a�$N;��j�������>ݕ��U�^O���͌��ɭٝ;������D��������ڎ���o��t�:i��Gء����6VZ T-���:8:z������ēsE��<��eʩ�����%H���������#�R"�M��/n�F	4X�x���K
g���׫���O����&K��B��^�s�­����+H������_	?�%�����Ks�9���h{m�cy38ގDｯ�A�Av�ť��\��Z��u����l̓oJȃ��A#p� 7��ÚO�Щq���w�t�K;�L{��SɎ��?�g<R�[K�BKȯ�~Î�۞�-С�H���1%d���/�s~�$�l����؎��o��Y�E�����n�����6"D�h4���.��]N=N�<'X�݆K�:L��Q+_�y�3�P/����w�h�:v���ӧ�ӎ�����i�=&txh�����ml��W�,M�ȏ�U���늲��Ѯ�ǁ��� �竑-C�-����ߡ��6���������hY|���(j Sk�d���E�z
�K3�$;J�Y�V�z�*->�=�c<9�e���r��簜�h���K�Y��C��B���\>�&�\��< -�PT�����<�x:*t(딁:���j��ў����%#�X��։�0��DP� ��������#�'�wU�t�4�氎�i� a��q����������ثz�Q]7?���u$P�Wj�(Z���痘P����TH�l�:�&���J@�R1�7�n���j0h=�S@�����d��z(����U�R
�y���ڦ����E3؉7��.�.��wn*� �A����}���&R�(�:�46��ߐ�@�w��_�\�a���QǃV?��oLe�+��\���������dh\R׾���%�v�(}��㬁�띴�p�T;����/�PW>�咵�<�k�E_�5Ȭ͏�������sN���8��`p�W �V�$n$��i�ʹ��@^0�2��K��d:&{>'����ek�F�v����u7�~w ���L�/Z�݈��������7�(���`>�~0�Ad����tդ��׫ʁ&����9@�
�B�y�yvnf$d�ƿ͟u��cE�s�M,h%���K�a�n�N�e��n��ߝ�-8(UȈɉ����ܩK0�n���kd���߯������3 Ll/Rm���y�ٶd$=�0�q��P8�@.֙"�f�|��PP�uE��pwioz�_hE1�66�>�"L*�=�x�i4�\�~�X�n6����G�� �8_S��� c6���t)�N�c� C��
�m<��t�tI���<u�G�&c���$4��\��ᶮ-駺���P8��"W-��g$�qX���á`:?�f�/LVY�,_�f2y���jQ�U����7��T5���J��B��v\(lu��jQ�O�Z�\a�z�T?w%j��J=��f���x�KJ���� ��G��� N�/��
;�0iEs������61��Cz��}bt	9�x�Q���/X������VS�Ww^M��1_u<%o.u�X��-�߆����jx��"-�S�dlk�$�'�W������8q�XϷY������'����aՂ���XjB���<����g��?��n�c%�Xy�/�i}wDxyYr'�P.M]A#��\m�`�����0y�	��.�?�C�5�����䢭��"�7��g[!
���_�S�DM�
�Zt�#�־�(K����$Q��!�6���Q�X�q��,ǻDU�B`�F8t�`;���S�e0�kA��_Ք�|��pA�LiO��H���
���W�Sk����ԅ��=Za1%����*rſ�H���e���ƕ�X��e�SR�L?le ~i�Y�����2.@������%�*b�k�*e�)m���{�R�~�A���<pi��������D�+V�2(��_��&Em&�����~��$Z��	E=.�{*�T^eV�����<�����΢Z�+}W��ĺV������:ڹ�tj��T|�nYO�=�و˘�![)��״7%M^=�k%6ޭ3Y_����pj�7�Qe5�?��^�8����c2����P�գp!�%YA"���*�\l���.�g�4I�4�z}�#��+{5�&�_���3�����W\P`���@`�F�8��i�Z(��!��am$����K�ӡ9Y)V�t���,Ю�Ui�"����ʣ��$�����砷��&�6U����H͡xMm�a����0���s/�j�l}jŶ�rr_�;"�yvV�'-C�{K2�G��	�	��V�V����Z�␐ �������/0h����߸��j���i��K�s��?�+fU�,�t=�����&�;2[j҆��av��
����Ɵ�v���+����;��X8���X��j��A~Yϕ��26q!���ml��=`�W{��qe��K�N��.���7�]7	��~YK7����Ԅ1[i:�ߕ��'
��?j�����)�K������g
+�H3{�P�Yb�V�׶�v��" ��B�$�"�!����|&��T�E��*e�M�{t<<E鯞�he2WV������f��Oygs�5a�P�q\[�w��>R3���w��8^�3�0p���t��K��K������$��2�j{�����)Tp�JE��s��jC>�'��\m�{Yh�#�B%�}�>!���-S��aa�	Y��$�$`���X��3
��8Y���mӿ�_}<��ƚ����u��_=���V�=rZӓ$��~���O�J[����I�Ƞ��b�!ũ�����{��;��&�}щ|�e�<�[�&��rz���ְ�Z�'ȇ��?���v�l�u<�n�	 ٚ�˓�"*N~v��c9)���J�^A�Dؖ6�	!kt>��`���E5�F�2��Q�k��:y�-���SJ6m��>����#�ʈ%]bo�O��n''�V�����;zI%�:��	bܾW���o�� u��!{���i?�<㕽��&S^��<ջ�X��,Z'�j�ĝ�~���{��D��8�-Ћ�:���Ӹ���>�wf~��Ҋ�a��l��a�@��k�irM8�{�W䁷L3��T��몒��D����{(���	���n��^�~��ԫ�{�@�Uś����	'p ���K������5����J������|�ũ�� ��[L�/�˳_,���/ݣ8�;��l�lQ�rRz�?�N�����L��|8<��1���`�R-a�DR����"g�G�jժ������(5�n�oj�,Pz�-���K����{?�<By'O�M|�J��TA��ؿo�O�F���;e��ўk��6��Z6�����|k��G�1٠E��A��j4(&i|���Pͱ=��h������b4WB*��3�b�wj����Yc�|���MӼ�4����KM<��F5��>������C��*�/w<0� ca�>��t?�e��\͎�6S}�I��'�]F?�k�����خ*SR��v9jZ{7�u���\�ZL����]Ĉ�0\�#g���@�1.�x�x��\��:|�u�8j%�C���%_}�7'	��a���5�B[�a�s�����tA�e���m��R���Q���I]=���UM���|�ѢB��GNE�&�����򦺈�G���V3�++'�R��-z�
݆�h�r�y�������]��4�	��|�i��aC�\Wa�䍀�
��K[�fiݻi�aG��
m�F޾�3�ds��X!h�do���ɉp��.��A����&@�=4�Q��'"¬����t�W��fcp�w�%MA��������M���.��/�B�m5�M�i���?���;�
��I�?�D��� ��'�
��?s�F��@-� 7����U�������p�*E�houVS�j��S{k��xٍ�
��ߑ �<	L��&��r�_	���݆x� ��8l�\K�����`܈<�����[�A��t\��(��P)LyT���DF@�aZP�F������b�Ͽt����Ù��B�}B��v��,s�n��vv�9+����ٯP�(�t��,"f������W���>͕�bn�mx�2.&|Q��K��6�(��퀮�n��i�\�y}�KdÓ�Ìw�e�4��y��'��o����fZ�w�sS��y��ob#�qgDO��i��hZ��+�lN��vш"��ȆQ�36�b�?Ʈ*.��k�-RJHK�t���C7��CwH*�tw�t���t �0C7|��s�����̞߻�^�<k����q0���̫>��H��������<�'�˾&���������T
�2�Lquo����z�Ur�vƜ�W+	�u%׾�3�*�3���:�+��:��Æ���u:+k�7�@�L�-O�q}Z�-�C�}�#�W�QT��Su�j7��0�{ݣ��6�ڜi�v_��@7n��o��_q�w�an{`���J8�UBw��on<H�^]֥���Y�iU<���^����G�d��>0~��ڃ0�����6�h�s﵁���/��I�֫Ω�l�s�X�@�L�6]zm#����ū��i볞��!!���P�:���5����Qt?���K"*#gE���T�(��B`�ѯ��υ����?���%e�3w��Sy&���m&�&\,#��~ц�u5�u[6�]��eR��<������u�ְt��FP�&���omOI��XN��&��|�tg�_�!_S���ϕ~��hRc��Xث��9��L�9�=Rl�� �~}9�n�_-�zb�AqV4��O ��N$^Xa���j�C�����wnK;f_w�;�7�rt�lodK��@yR������q����r{�uL��HE���5e�9����G�:�%�O_�ԤSS�v�U�D|rd�M�]�v��
9t ��{��K�iFՋ]?O�I)H_-�#ވIPe"E�O�����c�����W��.�P`��9��z}	�u#?����.x�J*lq���<;@Lw�wǣ&�] tI�~��(zN�l@�$d}~wj�R����~��(�t�<6�h�o��f�����#�v�_��ߨ$o�Ӵ��zU*ӡ��D����ץ��+\2=F��߯��}�82z���\j�1e}|Zs�~����B�����rѣC�zcF<��nEq�����RD�����CpX����v���/8�v�����sϓ$����6$9:�ϴ��M�B5c�g˒f�n���p������w��W�� �?���z���ew�`�F�P�1��Dx�q��z�hms#�
t�I�[��]���w��lIeBCrf�����Z�S���3,���۩f#9ٯ�p���0@��~d@�j���Jz��J�"Iy_K3���"��� @��ͥ����E�ʹ��z�)�n�8���uP{�%�	d�����v��ք�Xye ԕ%kAO�Vi���.���g�RF$��O��Ol^}��9J鸺�5�g���-��i�h��,�W���b��ӊU
��.�i�,/�}h*�����]L��v�7$�
sK\���P��K�yΠ� ��7�ٗ�8���X�n��Kݮ��q���(���V��M��>�Al��q�����������>K��*/�r�^�-ގ�1��gA�v��o,�!W�̚�/�N���O�}K5��x'02*�/�n� &�{4W��Վ"�O�Ұۈ�f�e�1�k�n�_3����W\8�+�ɘ��9�/��R�q�d�mڿw^�f���$�K�~NN+�~��_kE�sX�ӣ��}�����ٴe�ʛJS��Vſ�o�`������ Ԑ�0������$%�>΂w�96S���ׇ``�{7+~ؒ����-E��G-G�w,q�bUH���n��	�wf|�]��Q+�]�,�EK����xGE8s+*��ƴ�b�Q�|Z\5o�s��ܳTt�#������\�|Ͷl����(��(>�L�e��9�C��q���y�<�I2����~�O6�� ����VO�{�
M>!�fN�Fzh/�ߏX���&��m����(�8�|��'�X�eQ���1J�����W�Y�����͍�x���-�&������7���9�Hr.�������y֝�ݾ������0����-4,<�I�)�����4"��I�q#��B�&�>;�q_)�/8}�����Wu�wg5����)�)��>r�c�jW�]���+[u�k�D?P�x�m(�n$Ke�8?<��1��C�B*�|8�A����6=�Z�S !�o
��(�K�Пx|�]��st�m.o�m]�?\���d�A�m�u���K��r�pl��zFچ[׻-�]wEH3GĈ$Z��Fg+�3Z�VE�4[��|�~"�U����4J+�t��w�t]x�낢��<J�n{�x�ޥ���MS�7|!4m��D��ᦣ�l�����Լwm
���k�%y�.����4�����]�@��
�����d ��<���Ā-��Jo/;��S��R����C�DR�6�Le{��h�Ӿ2�jodv�'S.!/�K~)i�c���N��C�z��Pʅ�*�F���g�L��A�km�Y��v����Q %&�*��1�_��^ƹ�K�����Mf�Y��>Z'��R^��2���z�h����9�8��=:F��6�M�� `��Q~v��d*��Z������"{{�kM�'_C��W�~�t.�u�-��#,�/���ױ�ն�F�V�*������b k�,��$	�<�SV���~Z����h��B^$H��ҙ��K�!�C��l�
S?͜N���0g��}>���ƃ."|�b�a�c`̣�E��i�P=�[O}y,�v��}�z��9)��Nq	Ϧ�|����Zi�ɗ��Tf�9S��z;C��v�mch�zOj��SL��ؔ}�`�g�ƮE�ٷ��W��^�i�*���}=��I�!���E�.ٷ�Œ�2���EJ�}_0�}Ŵ�"B�EN����I0&d&��I�s�3
�9$�sl��
r��%���ٷ�u��7��1��P�����
_�+���=asw7��o,���@^��i��|�k���39V����S=K0��,��Կ�)Tnw���S�+�e��X��x����K7`F�n|�ɧ<8Z/S���[��i��ɿc�"V��� ���}<�a}[���϶�L��?r����n����S���Ŝ �<�� ���<O.Z<cT���L���m�[wD�e
$g�t[���B�,4�2ϋ��B������`��PK�K��
�So��>���O�F�J6I�1�:�޴�Ӽ!ɫLb�Z���VuSW/?�H��Ӷl���1��ɻK� ���p���
�����ڃ���'���y��ƘUܷ�������ʷ��u2 H���&-��\j��?���N�q��N��Xs�/w���m��c$�)hl=�@+�z�k�:h��w�	���f��68W�u��(�	2��AZF��^e w�<�/����g(2q��t�Y�K� WC�k��Z��+���eN61eٖ D�$Q���2����G�G8R}� >.m��ov�eɮ-U���b*��k���iKl�$o�.�hL,��=��J���q}{���[�\_o%���BNve"���Dw�;ۈ�J���s����+��gs
�Pk��_�h5�fȻ�"�;�VFx6��g���n"�$��| {��&S+NJ[�Ԅ3� F��p��,�\P_n��ٴ������:ΛE�82g�8�?M&g#z�W�.�LR�8�c#X�D�b�m�S���V��lQđ�-�M^�~̃����c��&�Ζ�!�frw����]I���a��:�%���T�dWVͥ.&!��2�ߦN�u'�w����Q!bZ>���[��h��6&��gFP�-��7#�`�ۺI3M'A�ﯰ%���ك��X��HIϗ��b�/��v�.qىnQ�w�:�Ӝhʾ��A���Mx���Oe4�� ԗ�k_4A��'�π�D�ߑ3f�����|�	��8�J�*�����O���6>}�Ѽ�?��dj����<���R���¡QX��PG�;{�8��-Mώ��l,τ[̳(}J�X�����Ot��C�a��kÃ�᰻��8�O�Cm�ȩ�:�����������E��r���k����&F�&��=e���4|۫o�v�¥���_G!�c�)��--����d���\z$�E��p''�}O|���(�p7e�>p�46����Ά��K)�<�j���e�e�1^���6
O��r�����\j���}-���XN��bES79�Yc�I�wp?���]��by�y�(�J�u��p4�:V�n	�vr[:$��4�Ğ���������2�J�u��GX�WAnTT�$����C�Z��Y�^��C=�B�F;B�:��I�-���˄'r3��-(!����vG��G�
�'���9��C��"�b���'�@7�T)������_7�$�R�M4���i���8��A�����~��x�5���LGyrr���¿��ǒ����2�������b�655i��2��"SS�i�y<s���9I��� ]�?�C��}�܋54t4~�G���=w<
���$	�	���J�u ��Gl�U������$�k�÷�3��3�$�`�?p3��r|v���ˬ@��ZmT���C��7�P�|��u�tY����H,779�,%�+�g͔�k�r�je[{�0�>�xhBU��?7���׷��s�[Yj�P=�[����~ˌ���u����#�k�-!-����f���~�ي����՞�*�112f����WZJ6n�j����=��� ��wj���#���YB�ӏ�'f-�<L�϶�ͯ�3�2u�)j�:B#���e�v��
@2��h���p�m窬��Y�s���.��P��E�__�����r%Ʊ6���`'���k�ث�;w��BP�ki�0���|躽�N,0��Ե�K��.���eU�m�ش'�啱�zzu�<Bh%Ւ^�ur��K��B��KYd�F-�Mu8�LšC �^�tel�A��fx>��(�Re����GP{Gd�8p|�c����lkS��0G��)�,���F~�<<�<p@������i� �Y����}��ۨ�=���Ϯa��ŵu��a����e�"#����e��Z{	��Q����C?��ă�f���d߄3�?�X��� �v�m�s���?:�73eeMNt-R6�^�I��2wgCå���g���9�?����ׅ�p��1m�\�*�̷�q�.��H�n`=��`�xR)�?��+2h5~x�M_�_���=���s�ۆ��'��<$�|>P�H�`ӥtok��}mP�t��b��[qj ~���Т�a?�0$l��=�=|B��|��*S���|����&v ⢦k8tt���x����OJ�o����`�O«��M���Y{y�F>1�(�g�Hxh�Ǡ��,���>�ؓ��ɋ�_�=���S�֮<����:��u��)>r{q��{��8�� �{<��?�mppO�(�pobH����+��9�>�J��n酭�[(H�o>k	3pl5�%�gU)��k�I�����bs����޵�zm��$�-UM2jɄ�/﹧KJK�n�hf��8f�N704��v8��h�T?�\����[���@t�1��6.���Xக'�!�@���9�N��9��N�I]�P����[<&|t���]�a�����h�_E竼��Uv򚙓o����~-Z�K���]s["�Ɵ�����Q{�5gr�y�M>�����C��!sv��
rQ�R��"v���A@J,?b�n�F��������y�S8,���0}��LP�h4���'�Y,3��م�ث�N���v}�w�7>-��xR��lPg�/.�N��D�F8��~����T/Q��u��{���OϠ���e$I�s)T��'{fU�� �H�[\�-�.b���h"z��j�c)���T>���G�t�4]�1�jbp��n��w���T���=+G)P4�O�>�[�w:�}e~��rZ�G%y����o
�]����*~�سԷ���Yv�68��hQ�����G���5�.������k"B�����fcawB�t���*h��,���ಲg�_\��ad��&/��|	 �Hg�����=l@�zY�j�x��[�d��l�l�ء�V'v�u��d���,~u��
���B��YTxͮNa>�YLp4���ehM|��lE�
z�־�H�w��;E��ڐ�x��p���ts��Q�R�[ܮ�B��N%���{E��БaJ*�>$	EE���d:���y'�=Ќ�EC�����HWٓH�zq����N���k#��4�<T�aK�*��y�uƏ5� �Ϣ���n��,��YUG�W�7�����M�ڱګ �>Eq����K�zQ0r��w�aq���\K���C�ʣC������������+|�~G�v��<�;��L$�.�Gk�喕��C\�Z��0�ϋ��W�4��k�7��l:+�����ʁ����O�|�hO��v�^����+�R����.NV�6�Q-�I,� �|����H5c�$>W?<����A\_��S�Ő]��V[p7h��������u�ު|�ý��	���_���#XEĭQ�~��4{ݜ��w�M/#WK���f��h��L�Dv4�6jp�G�u�ց�1���mOۿVsq�h��Ϳ����=���b�0;��}�a%��<}=ѵ�pA<����q`2(�4�lc����K���Ӎ �K�ր���S�~��\
w�45���x�_�9��yM"���~�B�+76<�|����_֓0�Ҁ��aO���u�Q6��λe}��Cks�)��j�-�G�~݋�ج���#����S��&t.0�S�wƖ���*�q���@��5�����k
�c�dW���,�?���)���Dw����ȃ��}kV��(��)��g,�H��X'�I.���w=��������]H5;9繚��R��s2�-m3�I}ή��u�ɠS_P�%&|�P��;7��d�MH��G:�������_d&�{�9G�fh�ʠ�2 ��$��M[CzW��js�vL���6J`� Z��}vo����@3��S.rh��'���y�x�	u���y�i%�ۭ ѢM|�w�����A���ǼW~T��E�1�8�H�V"��vw1�F�ʛa��l9�7������8ޞ����<$~��V��������ZԪ�'���2Xqkz��?����Q�HՄмH��҂��^~;7�]^��';�`'��?��0���O椇<JD���6��D���(֊���n��	�"��뵘��V����zޏ�0?�w����~�����ʡ����S0�s���ZB�4ʧ�(�a�g(�F;>+'$�=~�uX�9��F�����'ó�fnu�����'�A�>�,EHsזB7�7���8��S'/��:{B)<)(�f�t��xs�9��|*���ߪ��òh �����ё��3��7���,x�J��vy����,��#fKٷ�J���0s��{���iO�Ό����p� ό���\i|}�0����y�ѰiiWl��G���﷭FB"OVW�}�Y|�Z �۫!0!$^��+k)��r�ӳ{��cJj}eYц񏟦�ȹe���L,v�q��%�%V0��{m̽o�,-sN0Z��`����/(Eُ0
b��"�{��O���� r���q8�0�G��ShA��U��� ~_o�i���a�p�z������A� ��0Q����w@�-#�N]�Ï@������Y��5u�|W��,^�P�ʌ�? x��t޹�A@#�s�h�]�J���݃��%[à�4'7O�]�1��7���1LFS�y@�r ��HJJ��
�H]��`U4lGz]��v-�9�#GK �Yĥ�NfeEy�����	�r���`ۅ�g|��#���������z6�뺷������d�L�0)D_K-�H��/�z���`�EW�|�ba�Q�1��{�&����bCHxc3lp�3�\�s=���L�x!�+��'�^�@�X��Wɀ��������O!�Ō�W�MYFБn�y���k�|�[1"���:���x��Hӥ��m��S�y�2Z��^�U��-�|�qj� ����秬 ���ֱ!��q�(s�	8�3�$i��E�M����`�&tL+!��`-���[{�n��e�mV�Q����7��Q��N�?q�Ň��dzj@&�ĵr ח}����5&�o�	uVخ����ןD.r�m�Qte �YFv����o�OA��X�����"�	�/$�{��'�S�:9�l�X ��]��R]'^��R������I�x� ��Y��X��3�璂z|_0�� �+�ִ�Ƈ��O�(T�����D�=�ӹ�T�\��+S�4��낇h�)	�ɸ��߂lF������y8��c���u��}h����Z�E���Ce��?�/^��p�J�ï%��d���U����o(Y^4�o���G��
��z�u֫8�YV���0�a�X���t�T�n��Ͱ��aEY[�U���@�n`c'��Ç�o��H�e�ݧ(�%b�:T���Z��l�G�&W�p��!�,E�a�;�^���O*�l-�߼;��&��e�.D~�x�
�qYh+	|�S�뎹�$�4�j�o����5@�F��9�x"$@U���,�w��􌌈gw�ۻ���?�ɿ�b�?���f)�A潾f���%ޣ���+�Kڅ�Fo�r�B�m�?q&Y��͞w�=
�(;�Z�l�
knD���7��f�EvK��pӠ�?v��\4��T�����/*���h�����  Ѿ�|���{��#;�)^%~���gd�=���ǃ��/f�p�:�e�l����:3K��G�)�3�3D]�[m��cԧ�-;�*=���)�ge^����l��Ț`WW���9�L����w��M�� O�j���%l6�b_P��
��v�Tr���?�r�5������g���%Y�
���y]4#��toL�24�XK�c�i$ë��]�͞�0�c������j�)�-��Ih�n�ϫv�2���w����aے����2]�2��������*QAy�5-u�;��n�|ܖH���5���Ӑ��yΟ��Ͼ����Jn_#;j��,���ۘxĜ�>?�9����2pK����)��4hn�^�����6��kg硲����/�5��u�䭽�x��5�fm/��*Kz֝P�2�T�^/))F'np�7F'�9����E���Fv��(\�)�W=��0ɽ�_����p�3���ƪx��ӘhΠ�k������t�oilodd?%dtŔ�0tv@	��LXݧ$ߡ�Uzt�F�����W��2�_�:!#���sKO��s��&M��D� ����n��71�IlCB��]��X��� |Պl����^��L���15��\6$��19UA�����V&Z����)� e���TaW��s���z���>����wB"��GB��'M�g�*��i�Ԥ|�ܕ,M=G�^��۳&\�TrK�t}��J�$�^'�NB/��j��i3I�ɡQx��xr�[lT^U����/~s���g=���M��8���_�6�Y^�ӊ�����mLs���w�"U�S�Qkej�yJ�h	�A%�A��N��ӿ��Z��D��e�Wo?�7�n�s��@���(``�^��E�V����HO��M���!����s@���a�����y�����������ma�� aC��3�A��0$!�u~��L�yV�%k��S����l:r�ܝo���sݏl��Ч�[��a_�9��}�^�g�A�'�&�%�H�m����JuN��ԇ�O�Bhg����P:V!��<�z�|T%�2U�ͺ8�����s��L޺ާ^���;�ɼ�����ZgMH��"�z�2����g�x#@�QoF���_H�Λ�:\V�E�~��YDc[.�h ���:���β��@5�آf��$�_��vD{ܭC��{>9�x�)a��������浝�gMor��š��)�n+�
�b�c�w���Hg��ǖ�pJ]��YM�K�l���½�����Ό�"�2�����]c�I��9�o�&��~s��QN�v���V����e��r.���� j�EM�A���_����r�Fg/���O����f�(rw�*h˳yۿu��q�\�?=��Ռ��\@��;�5j��q�O��@:��zV{	~��\��,dR��A���W�/K��Ҡ�k�c�ɻø%����/?��3�Cgg[#R�U�GGla�׍��I��k�a93(�y/��pr���MK��FR),������xy?���Ɠy9������pR�-RPik����*AU�k�M�=3ȃ�����,���L��'݌�
�#&k�>fm�~Ye���C_����r�w	�!/�l�u�}e����t�v�{�-�"��+�^��Y��MR_cg�E��6����m���
���i?d���B��`���K�b��ii�_9���J�oy�k��S�8P���.I
n\Rvx���z��T�f�O��я〻kIF����>��PJ���+gp��k��҅���k��+���x���q�r'2��5P5�$2ƿ8Ch�9W�?ԮXZ��ɔ����~<v�=҅x����p��2n�nst��o
${壆5�#����d��2*PcP9N�[E�j��3�X��#�J�Å���2��R?8�=�N�-4���#Ŧ<z�=���ݙ,4\�5Q�.������L�&���p�,Hvx�X��t9�����������[�%��e{�X���}��FH^H����Q��������KI��gۢKl�0E�����Ժ`X~"�9�Ď���,U٭^_����ɭ�wi���M]������5�{�mT��csGէ���n�~���>� b��#3�y�d��_be Ǔ���~��� 8_i>٘��"��l�;ف��SH����Y�OM����*/���z�!�g���xO*�^�X>�Yd�(-,��`n�����	</�QհI�|I?�wJi�Μy���I4�@B*�~��SKn>��At��rQ���lG�*��#��/Ov�tN���m7&���4�d]��>e�Xi,tp<�/>8�vv7����-���X�&\p� e��n?#+P�ǪO��5����70���3J�;/0^l)x%7��R��r�a��+���:��-7u�ʧDH�+)�_���0�1��XwBs�݂}/�ָ�:�e�(���T�J
 X}�:��6�j�75T�|��Q͙q�1��Co|J�`n'�l;n���GO��uۉy�O��m�LT�]���A"&C,�m�{��l�6_���V;���1��R�m��M��\�@+�o3���9Ц���e�'���s �Y(#����IOEF���.έٕ�griV�|=��۸��gy��ul=��2��5�Hɭ�L���j��F��N�uM�Q���"���h�����XCI�y��t�o����=�Ñ�\;~`�7^TQ�k�SLeisG �z���|ઑ-U`Ż��~��-1�E�BTʂ����"�Ci��3eI =�8"i�4j��乺�V���~�_��w�P�|�%9I������􇭀>M�*yKKƋ\�{����R�E�#H�p��3~�,���&�0��������X�)�#�W���s��Vk}c 0�>��߁�Mo���P��j��`��n������Q�����#��ە��y�o�B��i��7z���4-�G�-�J��H+�����9�K�5�E/	>��c|m���Zǯ	~u�9<&��$�!s^�L����Xx�"��e�̴LYl���,u�y����xb�]hT��G��8X[�k���k��\��}�;�� ���Ll�cprUp�h	�ݲ�ȅ�9k��OA�~�м)�LD�V .��i����j��i[p�#�/w=��7�,HS5c1�hcR�?C��%�7DE� q�u}BX��}Ӵ�3{1�pji�mh�:�0g�u ����Ⱥ�tvjy?��_޹�C�q�� t�������ol0���ۛ�x�:��qu�^W$�4�[���q�(禅v ?�7F����fkD�5[{�c]O���H���O��WN�x�s�\k�Ἰ�'����,T*������O�����f��v�:���Z��ڮH����� W4C�Y��T��p.9U\���)�ť����=��|>� ����_������}F)�'?��ݓ9(����b����a3
I����'?�#�u��֥��8��>�㿝222\������,��!�W-S{t����ii�j�̀��a�F�ď���r�@H��y�����Քj�mc'<sc6�`R��fq��XG���F=�M�9݂�*�f��3mWgS�4�ȋ�R1�O�#�4ٌ���X�����^w�.ه,F����?7B2,����v��m�!ُ"t~(!i-�W�����%�T��};"˽�4���1(����-/~���&�f�tF����FKc^X�{E���M��֌���'QQ��$R��^�ɸ�_rēw�||�tF���DK�c�DE"mL��BvD�A-ˤ���*K����L�#l!�r�b��g�����*��G,�˨-��X�FW.l�����J��r�}i��u/\\G�		��@���g��v�����R1�������,�U&4t�ڢ�Ia:�������ٕB�U�"�&疢^@r����D�>��{/SXC(�nبS�Z+E�\�oI�������^cdi1j�~y�PSSg�V�2擓[�����u��߫n-$nXYy�tzD�2 QS}����Ǚ�����!9sIa��U'����E���*���x��W��4'��g
�v"����	�R��g�Β�w^,gs��I��"�]e8���b�����%�z��9��e|� ��B����_��-�;����1��޳�?ޚ�Z����(}(�M����0Hhsz�4y#����h��-���l���޾�E%/���w?�F?-�Ol��-AmC�4�I��}�t��ħR8!���d�,a$�����I��������<v�b�V\>���/�p7J�K��T�`�������oY��WS��X
QZ�lI�W=I��I��zR��i�E�n�Ɨ ��>Hb�pB*[oE�,��@���>��k��{Xfm��_A�+�qn�S�����[�J�Y>�nqF�Ҁmc��U�/�W�X��D�fp�qin�7;`�����p�>��8=_̵:�G��,=��Zd�Ǔ��A�J���02ob"�A��Y/x���T}�ӿ��*���,�a�����A�0�@A�bb.���`����)������6��7�z�
�ysU�ӝ����)ɊU�fT|��=h�m�=��x�.(�q�|?=#D���JrtY�M�I�2%3s�Bcz��E�O9%��:��5��$߅�ji$z������2�V�j��v�����/�xm�OƉ�"
��= �-�+�\�)�o��)�Z��#8BML�z��J�˙��U��V���y4-=��(�>��BF6D؀�>u�;����S�]�6�H���]�teJ°��m�PfO�3W�=�� �J��x�Ә[Uە>�2��Lr��2��B�����=r���&m�R����4��z�G�OvM��p(SѸ(����T���lxvzG�{,�!­�7�"q��X����sEֵ{��O��#�P�
����r�^h�yG�(�֔��9��7�椖c��[�/i� u�����I�@��څ��
�ͦ����b�H�~\;���r���Fk܉�ꗈ-��	���hc��$E�J�qD �����:�g�zQ�|
��S�����<�OCⷛ���G�0w-M6��qp�0����5����������8:�z�����e�T�9a�܁$ �B�`6�G�o�:5,r����-)�ZY8&$q	>�B��t����ݳE�9�q]+�˚��z��1��7�֬muX?%ӝ�L�z���pH��{tm��kY��UIN�(³]�z�딅���f％}<5��s):6����K�B+�3���d������y��/����-�$�7o5����)}B�H����T3���OS�̑,��͓�c�Z��"��e��1������*�㬾a�cd���1���Rp�9�}�\���S�ʣ�b9PIq��ǟt2�W�ϡ?V�u��wo4����m��,�-��z&(��OM-��Me\��)s쇭����\Ə؍.��ɜ��Rl����i�s	�±���u I/f��f�C��m�ף�,�~ݏ1-�6��ds�k���W�4ρT
�s���/���~��ޕ������X�/��G�6=<�ձ�R��i2���=��lܒ�9�U���JQ�ͳ�M
/��޻F�^����H�7Q�N�ί��_����>M!<"x��������2~�ٶET4�x��W������a����WBnQ��*hB�ޙ�2j%��s�zL����Y�32�z�T�T�ͷ
,nܫFVxӿ�=�ˌ���l�R6�$h�Kv�'*��ڝ�^eT)�u��d"�����.�����O�jJ+쩙�*Fl=�<��o?]�z��^��yH(��
7����G�맄~B��v�LDg��-�'x�C��:_naCp�.�/�dy�~�Vn3���,d��e�6lk ~S��,we��(kP}~E:G��܁
TC'+\<�K��$�+��_�!U��W��+C�M^Q��Us=�W[+��߅?�%��d1�3�PO��R����7X��1��L����԰�d�z����l��v��ϑ+��� ��2UN����۫&Q�2�=�9	uE��]"QnR��4��
��d��rs+�-�E������z����N�5�xz��MaZ/V�P
a��-0)"���Qu'��+3�8��~ ցm��yy�i��P�sm-y�D�V_�#t� ��33|���z�r�x�9nw�v� Y�R������el�����1����X�2؈ϧ��N.�U����N��	B
�>Pð�<ENW��/ƨ��'�vu�{���ϫC�'Z4�H�kf�R�dH�Q��w��.�P��(\E�z�}�;��ĩ�^���ux�ڦ�O9x�s��	���c�����'��֢�e>�-���I>,�UP�}�$������
��D "��'�L�El���e$o{��13q}��/ �O
;1XwKM]m<� Nj��^?yg8%%�V���[�Tb��Ke��x�/_�sd6�@�\�3�A�N�ϐ9��m)��#8p���	���MAB]7��<�i���;k^��ZA����/��g�o{_ �����c|���{-��j5���OP6%��4z0�{�F������0��}�L$��<��ڭ-.��F̹��}�^���<ң�xJ��_'E��e��݁�>>�Y#�{.�(���)#iP#��9X(��6�e�����J�����W@G��
'V�w�J��d Z)������E�+-5q��<}��~?`LMe�B���	:�b6녳����8��J'��a"&��\L��ݹ�r�484�u{�1�F��.s<��jWt�g�$�����#-�2���g�0#OQߺ{:��l�y
�
��i�{�խ���2ѱ�[}�|^"f<﹞�4�PbF+~�<uȩ�_;����68�����B�	�f�ք����#K��k��8��v��r3 ����5��j����7��Ũoy�K�.rA1sܭ�(��[(`�Pf���W1��O� .%Y+�D��½��/S&��*��rV�&5R����^��x� fː/E�
sk`�ґ�+��.�c7~�0����#�N�I��f��ܴ���y�G���J�*x�����Q�����t��5�}ͭ�|B��e[��;���_�[k�'��bg�M}��7���y�B��Iٷ�]CY,�@ܭ�W �D�x�7r��O�h��[�5�=]���.���b��|�Zm;�gkm���iN�<,�O~`t<��$�t�qϼ�Nkp���:Ɯ�=8�������zYR�*�J�9�v+�к�v�{t�D6�w�;��Q2�isӷ�����:{sL����Gsؒ�q�ْm:.B��Ч$g/�M�hHF��&�a�x��We(xPV�M����j���y~���?Nٛb8n���ܾ�/�>%��M��kB
�C��}[n�P0��H��ga�� #��װ��l�m�[e$7�3)aA뽁��u���Q�*%L~��>
�
_�W�
�H�WoH�ƍ�)n0PH�9[�^�9�:H}���G(SJ�=����<��4��C��7Θ�Ǹ�<ǭ1�;�bW+�����^)6|����b��Fڿ_�u���6�)�n����R��	�O^����g��g}~��}q�ԝ���O��n��������hv��<�Ĵ�Az���~1��j�"�x}�[��Y)����%s��-	�AvW�Ff�r�QCX��G���%�ܷXa@�/��/�Wd�D����rX?�e��R.�J\CNZ`��.��&DAb�4�s���D��֎o��ZW�ؼ�ՉgC�k�}J��l�>n)c-�V��@9K5����nJ��ъM����س�����h�TY�c�y���.�jXf����@�h���Q;���l���$۲�*F�trA�b�/�[9�
j;�E��OiXR����
���Z����S�IN&	�Fw!5Y�"���[���k�	�	�	���݂����%��;www��w�C��}�}1�<kuwU�U���nM��j �V:�I��f�>0i�%�4�F{���m��_�?����]ߥ�WnהS>%|�%�G�ѝK%��/���<��!������y=�V�e�2��zu�U���O�ǧ�@�gW��@�����N&%#N�x�~'-w���ʋ<)ꍔ�9q�ӎN.E�&���$B9�η��׉��@4cJ��ys|Iv'����������y�jUT�]�8�G���#�u������W���W�|�S7��B�Ј��%z�D�EF #��$�q����K��@O�����K�h��}Y�?���W&s�CL��P�.��6YN��6y�"���n`V�մ���՝������][�o%�������gvH��݈H́��F��J�R���k�:<̱'�k�6�|�
���^_?�1F�V]�h�T�5��1XS��'`$��M�d��BX��=57�_х�Ԃ>��r2���՚�%�|�6�2�*Z526�҄�;�0�8(��5p�E�wG�������q�yW ͳAڑ�YY�n�
tp|�q�]`_��f���ߒ�� ���óI"֟Ύ�X>���/��.-�|3*�ߛ)�_`*ס�����9�3I6��0���h�yު|�{v���Q�o���h��м�FJ�TmX�]�y3*/J?IwZ6����-�qw���Y�B�7�y�a�@�Lm��_N
�������Y9�� T|��T��Χb\�'�`;�Y�>/�X�{�y��/�����蹘����!D���s��3�*��p�^�r�gﾅ���;�6�@���ᕁ�R0��b6w�=
w��wAAX2���^}_��ځ��±��.B�:�]X�$�lu1ۍ�%�7�8+��6Vx������
�g{�z'L�����i��2�d|�c���,+�>{�-A>�7p/g{!Z7�u���-�?��e!ѷ���sw���ɍ#ً��;oP��Ӎ3��B�W�pDC5�0��a�ydy��'I2�J�#�0�BFW%<�#F���,�R[ӕn�R�Ȳ�w�x�}���眣 jw��t΄��PHm���l�ee�7�Dt)��\(\�� ��/�hKX�"�m^�g0�z�����Qa�o�����ٸ�&}L���o��l���~fX�H,E@�p(|�8���C�)} �#.��l�<�행,�#77�c��E�����8�bU�Z��²
@V��큶Е�E��՗��~�b�S��fFhHG6^QC�c�
w����o����rԔ,�x�r/��
� Ys�r��T�r_N������}I��u��ز�j���S]�4NKӾ?��0�lI�+J�/�*�H#0W�6rҊ��l�����%Ue��ʣ��t1"�qA�{�£�wv>�h2Q4��3٤��@��K�o�%�*��Ue�_!������gG����2a�kț�@n��J׻���PGBe��%ue(o�^�V7P�jd�}p5����1�?_���G.(���>bx��96�����*�rme��,���;O�>l�¿�c��S	O�f�^�DFQ�@�1?�XZ��X��|8���b�7�v�y�ί�7������A
�[���Qc�J�&}y��@������v�z�O:���:g��z��u[�����3��T��`�����C�I�E��^��� ��x��E�"��[��K���)��nR���"ŝ�J@H�y�v�)0����1{��͊��>��̻Hg���������t_=8��4���|N�u+U��J&x�v[�z����Q���D���qb:�+e7_Z�����s�u���q�.�������j�:�$^�E02b-��˯^��*Z�|x�0PV5x���p��!E<�Δ�%̕b���a�޾���M�KZ��h����b�Μ�_3_{�Lh�wrM��ɿ�I����ҕM
ϭ����D��d(��0	J�&2���%2��V@�߹�J�4B�Z,m�s����}�����J�?n�Bv�v_��׏��[�/��f�ސ���`Y�(b����!�������^�%�M-�J-��tK]]+ ��p��e�#0p#�H����NO��(3�WLԲU��|VՓ�#0�3�ނN�,l������E ?���-gd@���l��I/�!�@�W��ZB����&'�e�t<�S�<�n��E�mݟ�h�{�&f	��_��j��l�j��n�,wr#&H�d���܃��1ݬ��E�Oh�û�?!�7����_D��=tW��8$ߪ&{D�i|NA�;�n�*$��^d��ĄC��9}���rC�+YH� ��ԭ�\}������("	.7U6��>��`��).�۵!���.�l#����$-c��b
y`t �ǏB@q����uR��3x��l��`xKh���V�F�Ջ�]Z�B�5-R�wX�X>�F$�Oi���Ys�D}��2��t �x"���.|y;v��0md�K&HH���i�a������s��,9�2�i\b���&�൅���WT��=�2b~���S~k���?���W$e���c!^Kx!+��1�22Ă��8�M�Q�i���]����õ�������~�_,�U�S5=SU�#��⻫�uM �~��8�3����ط얘���ɝG���NR��4�E��K��v*֌��o�����\:A���ȥ\��/�d@��MJn:GU�V0᾿/����Gd�бg�����.=����n'=I?�D�}�\���+e�D/ө#N,�)�l����K݊�~1�H�.B=��@����㍟�y���i�
��Ej?Sq�f��ęˑ�0���x�[!���������4�|���UxH2R�p�~�/<7���O�X��d��NU�P��4��p��L�R#T��0�:,|��g"�mc.�=#�x�!I�Kļ� t(
{�5Q	1Far�0{��Ts��^`x�c ��@�vWa���&ē�o卵�A�{=���/�/Uf�`�}�x��#I���RUm"h�>�l.n����f:	q��,=��˟[7|�HJ����
BOZF�Ֆc�|�m�IJ�Tl*!�G�K��ߴ��ӥ��It�2:o�Jz4�.��uQ�5�Ƿ��{�on�6	�j�)�6�:��a�SǷx#\@�7�����Zr�A�YYVu�6-��3VVvǚ?^M!S�y�nm}�t|��6G�!�7 .���AQv���k!<%��_-�^���g4Sh�����^lo�S� �g��F��p��0Hĝ�_^u�3��<�=^6O:A��	И1�Ǒzj�ׇ���S';�*�kyzNW�Z3��C�˾k����;|^i=&{�)Q�%�Ј����-,���]�$�ު�>�5$i�*�t6��άZ����&�x�o�K�ݹ�t�7�V{�Nh�]�4v��|�/P �Y��]s�OJB��ͧ�ϣ9�S	��	�R҈<��S�I�[�W��QLZ8ƭO���[n{�OfB�̃�$��N�]��q.�ۏa;�<�J�v��-hr���O��0 �ƞ��ﳶ�ޭ��w?�&�l��!������w�$�����IP�5��hT9���+�Z��p�o]U�H4P@��*� s�g�Eb4�sM:W��	
u��EL%��p��"W�f߼1O/Yo�X3|P|���W"�W`���5HG⺅���陲	�5�}Ǖ�� �Dyʴ�^;��tFxR��V�v�{F=R�\QB�N4r���֛*'�..)�d�Ƒ�D�
��޸l=?Vq(�c��������t%���N��ybe�*�q٫�5�8�4�]��xt��X_ˏ�!~�VBo��*������8^��Q�tg��)�b}�(�@7�t$���/o��"��.��:�ce���ȧ�w쵑;��XC���/͟��r'ύMLu�A�:u��5-����+�k6,�O�����Dr�"�C>�{ZQqya��������Sz1�X�t���=7�A��[�p�I���#�YY����l��]��;��O��;.ĪkÖ`2	�!��K�l�jݴ��'�8;⇌����-���ig�>��~A_�P�p���F����>+�@������¿��e�������_\��5p�c�
�m���b����a��B���Gp��ſw�Y�?�+�BQOp+�z��~��6h����?����v�q����%��.����:X.��N�G�܊�ഛ���B�s
��g0�jmz8lcFO�]�TP��g�v�T�����_i3&Ls=�=3tb������4��#�!W�j~�Z�L�`�P`���6/-l���>C��]�8`Z�����?�5��===M�<�GW�S��+�j��za��]���_�������=��q,��d3�����p�B]����%Md�\9�	�VR?�+�L�h5��}j������[>���B�D�aȟ:�P�ٞC�Y�_	JJ�*�_�:���V�jS*�edSXôm[���ሞ��*�ϔ�:%��9��:�n`|[/�@���l��KdH�9l�9{��<������L�� V1�ii�ߊ,���:�X�l��!|����Z"�&�x	�����f�^]����]"�vs��r�[o��=\Oʥ\$�^j^�E<�l�ݐ�>d����|����_~苵�c�X�l4�1զ�k�ս��dEW>��6g_}[<�����8o���L�uI�<(/w9�=��$��S�"K�$b�K������{�˽����Xo�s�)n�W6�x)�m�]¦��z���O9�H:��v��(:}B�#��;�:���:3�nZ�G� �T�T6`{�Xv�G�/��E���coH�p2V	��*)�
��1ȍ��q}+�u��7���ut�]s�]~E��r	��Y�o���Q׫K��}�Mk8?�M�Ŋ�� V�
�?��v�(z�ܬ�
������%6/]j�t�]�I���5x�R�.' �/��sz�疸i�3S$LL������w8�#�3԰�S�LUl������{�T�l�b�c�r�*c���>�r��&���6�sx^w�yg�����X��_n�&�����2�Ɩk�1���V;	t��/��u;�y^�u8-tjG���B1�ΐ�s�h���3�u%q��� ��Wb�Ƙ�л�q�e��T�;����[�է	�7����[�T��C�}}`�H�1{nI;�Y��)�Ϯ@��\������ٮ�|����o4ϗ� �a(��tG����͆7^f�8�y=��^ga� �tTsk�$ݪ8������ �J�� >�����G��+����C���'6�����4�n�<敐Bf��X���.>�-f�����uYXXe_����>Gو�L�/�
:x����D��v�����5�͏��s���s~O9��ɑ�NCFDz�!��"�B�mq��=��F�qW��m}���V��� (}"E��?4�y�\31娥["M�hӯ��N�H�KqO|�:ns�}cQi��?@�f�O�]\��N��hꈢ.Ǖ%��1�Œ1jW�F�Sc��Ub�jl��͂s�G��V�Z�����������uz��;!���G��f��"*}��ͥG�~�#hʊ���Q�U(T(1���s�aUUUy߮Fۮ��~8�Hj��g�y�x���W�{RѪ(���n����u1��I�NO3�ca�2��*ǆ�0��n�����o�8�{��:��,�OP��)7���T��(��\m�dݿ�
�Zٛ��M���V8�dD���HZ.��Xn8X0��;��rB������3ÿC���%'�����zO�
JY|�l{�R:تH�(p����)))yy�%U����)�OYQC��b�y���J�P��v3.B�������)$JEU�ִW���{ZY�*�����6dK�������ڪө
=�@��vN3Y�Lq��u����"���̝95uT�$�-=1m���k�P�t���?qx/{f`T��Z:<;1��%LL0ޞf�	~nXTC�gו����D�r0g+�~h8�Q�QS�QV@&�7���LJ#���P4�$d⠴2.�^��p*� ��ϫ�Ło7"�Ǩ5X��bu z+ &�}Y�+v���c�f��e+�����\Ԅ�� ��DaD@���� �N�Jb�=H�-S.�iQ%Zv����H�/�O!{�:���}Ucv!0�9:�u�>ܓ���F����Q5�z��`��|�]���t.TKnc��{/m�8,�4Ĵ����<;���!�[��٬n�S���X���X����@�{�֮=z�)4Hq����8iD��
����)�f�c~`(O��V������o��:�Cf�rR�(��CAJb��T%?c���+[�!�i@�F���Z���{+OK�K���r����j-�M	O%�����C��&a-/J�K,ȵ2���FN;�����h@�۾��vT��:5aA18�l\�p��w��AR�t�	ES�$�$��@Z�s:r>��7:$2����
#��4���~6�נ�ـ��meƅ-K~��ϮPR�bǄ����ňfi�@���FZ�'=���]�<[k�ߏ�C(�1�eo|Nv���K�7�|���i݌J���m�H݁i���o�q�g,Z#�����x��7�J�rX<e~���:|�Ƚ��J$��2VTLa=�3���*�(��=� R|�z��V��B��~߄��yo������Ə�v��OC�BQ��?E��,��2�@LG����{�/\�i\���"�.��m۳m'Ǭ/�1]�p�Z���~�Ȁ�f�Vٱ樓FE��3���@�UN��9Ikd�cI��:�_�w7�?�,�e+zc��9�b~�e���u�贡��i�_g��J��u)��A7���oƢ�`�h\���g�C�������saP�I��6|-܄d���g�\�aX� ѫ�&��7l�x��k,ȍ��j��l��i-C�`t<����]���۔q�IP&� q������roʑ�Q�xo���6k�	6���SZ�~�"����d� ً։`y���������pVcU�����WS���͇�֐2u�0���v����}�|ܴ��ifKK�g��Y�b�Zx�lq77������+
�-C�0�
����͜^��֝��AT4�13��R0�����	86%S��S���-��[��<��h�
2D΅0tӭ�z�p�8}��q0�b���Х�h}�B�'P'�Q!��8���(�m/ɑ�<=Bۨ?����v���\j�d"Ű�"3s�_��UQb�-���P��:�B[�2�h/��Ծ�M�o'���` s�k��z���>�	}.��,�o��(�����<۟2�]6V9ˣ�f�S�?�Q�9���2rw=4���@u!P;xb�������ɰR���|J܎x$z�׽ō��x�ȳ}��9�]��*�&YԔ��񈠉�37�ѕ�"����}D�����p9����{���jC���2��B�}�(�m@;�j��!ENZ�N,	�N-|tA�� Z��Zu��^W\�`�E��̣f�2�[��}>4c2Rh��\Q��亦{���=��83>��Q��͋c�	B�?�!���ՙ[J��=��b�8|���R�a�4���4��tF��Or��sҊ�pP��5ULN{��T�m۶��eF��{Ѳ�r�{�1�"�0ie�3�5-]B��Iеƍ�2������[�:���	����:�R��O�����Q�Q��DT�a�M6a0�Ｍ�п���:`u�o�� �v(���H�Whlfuܧ�	�S@YW��E��=��!�"��/�X��@ԭ�_>7��C�ĵ?�c�Zf��o�b߯R�[�UU�|��ڋ,!�N񳧉��+�δE���y�-ͮ6�(��LP4��oR?r���j�C��.*���Ɵ�����
ϔ��3�H�/���f\'����cL�cp醃�@|�vW��;E�7�����D����u�yx
>�H�Gx�$Xu��$A��Ny��>.��u���2�����䬓��fX&�Au�����Fo��gy��ajl��Q��#��������u���'��U����.�(���z#X/�'Ib�F���>��	�eC�'4��tZ*���߉�^����3����[�m#|���`f�>�	^cS�͈ʎ����u%%�:�K�0e1����wQi%���߉	�3��h�����
�щ�[\��o�ᎋ�U�O҇K\�Z4e+x"QB���c�^"a�޶uZ @<��*���r��N��c��?O�KZ�&9ݘ����:�>��q��f��p����v���m�M���S�1�m���W���`� ���,���zE1=0=be�����
��1��+!�<5��N��+��
��ԁ�T����Ao�*k�B���[�z���i�i��E#:���X�b�!8>~�deG�
�P�iD��8;�qO"\Wj�\����b����0��ϟ�5���8cD=��ao�jj�r�'"��A��p�j��ِ�i,���:���t���� &�DLC�6���n��y��2���ߓ'�3}]qF�*�HO	>����tA�k3��Y���5������p1<[���X�በk�M��y��P�y����"����)��i�ݦ�/^.���h�3�zn!y�׌)������\Ʊ��ت;a��oN��O��;~6�ۦ(�	�g`�����;�[E�u)�ܪ�����WQY��:q��=�=fnVe�B�Z!}��v,!@X���f��8���{i �n0V8>��U6vf�8��ﻍ,ז��б�����m��	ot���$|�ʎ�p�ynB�Ft��C=x���?B�ן�&�|��js/z�۽6��6�x5�/�Fͭ��x���8�[��9�R�I4��D���B�V�5�a��7/b��5�t#|-�17��6�ks�P��I�F��91���)��E<B����ۘ��2��6���8��đa�vW��K@J��o� I��������oΔ!�13xӋ�-�W���q�Z}�1�SR�?~��qi�q�x�Q�u{L W�47{.⣐�p��$T[�Q\E1L���n1e-;��  ���K��k�]�ީ=��CA��AJ�O�I<��)B 4n�-����4q,�v�'&!�l��k��u⑊f�i�>:�
�۪vX9�D��&���g_���&[�'�Ą�L�r��V��fi�G�AMĕ	��wa��ߊI*�S?zxbL�홸�lzņq쨭Ȃ?��� ���=�S(7���R���KzA�IC����,�n��[Z����&�����A���Y�R胱q'���?��K�\)O�����8��s.���S��i@�z��xs`�d���K��vR���]�<�i��e�c��ܤτ�L�zFc����d����~A�8�D9�����KZ�l7^XuW����{L���.�;:n"�x�3�������
=K\mޙw��2ԟ�{ �9up΍7'���ؼ��r���d� N���rI�p˩Z�#"�X�lGű�"���v�VRH/�T�<#���/�>��取匣�mx(в�օ/.�c�:�J�]����;���H��񋶜��4��������r�.�3��\�/Ң�4$�_#��3>rRH���+ ��W$ۓ �ׂ�5��~�\�Q�?����%�� ���Сz���f����9�;�A/���F�sW�A�P�#&ȱ�sByub���x���Ϸ66u�&����, �P��o��85�Nq�ҫ��`xf��
�{&��T^���W�s��Z�����!�ҧ:�eI]כ��|��\� �͓���i��H�	�&1;�E`wW�U�k���������ʤj?X���w�7��s¶kl Cc�����n���]�|������ʳ�g���5;V�7��Xn�ɑ�I0������8��+z���D����;y8��#�ņK��ai���7��,�r(Vp�c]\Һ�ߒ��"*��#eYӐG
>����𝲊ѹ'?9�y���I�r��`��bu��%g��}I>�����+;�����y&ܽ����P��wN߶i���۔���Kf��]X�5��uԒ�1����驍�%���h�N�]�Ѫg~ �R�e�ɡ�E�8�I:�AxkO��e�.[F��j��{W?%0�m�W,k�� (m�Ȟ����������y�=9�s8\���o�N�*"v����,o�>$�����yG�)�`)Sb����tS�t��rR�]@��$���y�����F:"o��"Y_o�֜�(�K�(&lD�iL�����hw������B�^�J�^V��Pm׋Nɯ��
�,��F�"���H�]1wN	�R �r�l�	�n��SY�F�<��я�N�M��Mf&��p]ǰ��l�P��I�c��kN{7c�z`�!��<�Ju���Qv�է��'���x��������*���F�s�,�BF�Om�r���c�V��c�iZ]*~�^���:�/|mŧ��;���{��/����ڝn��9,a-o%ϊ�
��_ȩ����8J[��-O��o����ȗ�ײ>n�=�5�m�ʾ��v` �ҋY�v�+A�~R�N��)EAv(j�J�����lc|��daw�� �ûKoh<�G�E�`OX��d&��ؙ�<Wܨ�9_tZMj+�p ���٥�u�S�D�V��Ns*�E}�!lF�����鉩�)�c��'�sTSc��5C8W�a&\kVn1�1�m-�e>/5����/�$��k/;N��:���v�@z�:v�_�+K�brk��	ܕ'�������[K��j����}�V��|`"Q�̄�Q^0�E��3���+*����lrvus��|���r�τ��h]P=|���ֺ�*��hv�}����bs4�&�5Xu�FK�y�4��]���t�r�NHNU|��G:�[K�PG�P׭�|p�����a:	��4V�Xᘮ�쪡���A��]��ݦD���g[��C���E�r�Eޛ���d���\���ߔZ�{SS�`,�3F�J	<$�k0*���)KUx���,�7���T�ї��ǖ���rw6��H�X���W9ǼS�	:$uӊ�����-wˑ�uq�����/,�z�� b�~̳��< QΦ��� a#�ު�AY�4M�c�ijGS��=���Iz���������k!����;�-@�`,7O�;��;*,u�˛�]�Vۢz/׉_k*!V!��	�>�Ih$�w�>����+T�f�P���bK�r�[ٱY���m���L�c#WY�h�y8H������O3��5��P�m���i.��q꜑��1�%�Cz*��f�st�ݼ���z�s�]-#����d�S����gh�v�oFx5�񃞆�mU诶�*nr?��k�.�O	0�*���C��-���d��*�ucK��ǜ~�u\���I�{����,ß	-?҂�x2,
����GL�w�E�^bE�	2�yBw^���O���p�樢��L�b[��V�֗��Q>��.7�a����!�f�		a��8GY?3Z;X�F�g�*=�wp�(�\�^]�6���Q��	�-������***hg�˧w��_E�ߣ��CK�8�V�x�퇕�NpӚ~�[J_�73TE�����������6�T���\B�GsN0�$Oo���֢XPk���	**6h�R�l$��ӻ|��񽢢��� �;�?=���aP�����b�gS��C�[Γ�'TK���+�p%s��"���7�Ǭ9�ܚ�Z6���z<�k���gJc'c�a�Uy�R9Ĕ
�
)�TD���>K퍏��Y\o���Dah���^߮P��Fx�ܣ S�E�=OOu~�TP�a�Ln+���H�~Q�yFME�a�۹O�!P���?"a���:�.�_��u}�i0�㨇*K�zSt��/g3>��&���=����K��$V�������v�r�4g����]v8���D$L�Jձz�6�H>R�]hA�E?�4������hw�� �'���cSk�W?�>e@J��U	D|Yu�c|%�ƣ)�QV#yTw�@^9�w�޺���Qk�����Ht}��&�x���BD���:b�XtCT�M$����,t+^�c}$��:��B6�%,�8Ә��j�z|�k�ۊ��uW����׀��)[x��)W��'��G2z�B�	;�s-���鱳���Έj��ВeA9����
y��_��K޵�kA�?n�r�����|�^�FFU�<D`%�_��6Pc����F�o����w���t�i~��LP�e0��_�堟Y�P�%t1j��GR�!�D�b�A��h�Ȁ��u'>6���%G�ng���U� ֆK�m2�r��<�`͟+��K���z��e��=ka/��
��T_%!F�]�=h�V��*�\�=���=�s�Α�����y&RM2~ .�˫��˼`oId�����������_óG��J�Ys�3�����Ӊ������?w�s�v����_���I�%�����}4C����SmM
��IL�-z,��C�;��K�4�yd!ǅ��Y/�=#F.����Ȑo������g���Κ������7#x��!7��NS��h�u�w#�#m�n�k��V��g���G��DƵbF�����lU��ӵN>`A��U�CUv�E�3F|p���mu��2��YB�ն�ۭE��d5Z�ؘI�����օ�b�(Hc�Qˆ�]_�	!�6�t����eLJd
��	o�2��TB��\[�C��+3����{\���r�c�z��j��g�n�3"Ʋ�5�Mc��ox���bJ���<Hx��z������Y��
�E��;ڦ@BA�_|��b��k��^���0�#'�fb��u5�F���B)�	!~��M�������_uOɻ���5���DT``�$G{FY��f��^:ua�����I���%�#�'�[iP��J"��00��᠎�U�K�������V���Y�3���=;L�Xl���pt{��* �T���'��4�Τ��� �+/��<�7^��,�n�:.)K47��a��Įe��ׁ�P�9]�W�5wۙ8���t�Z,��+�zv�w�N9�G����4���k��T0fͭ���L�ke��-w"���ȩ�\h�=�F�d��c\|h�D��klϏ�V�و2��/�����@�\�����������i}����������j�`�i��ϗ^wg#��QL�i�&���@�YY���f���Btl �{�5g:�^��D�#�lsfH��C5sW&��Z$£��O5�g�@F��k��cm6��$���yl�uw�z*A����`�SOm���o�7��NUX�>5_	9��c:�o��K䲓�"����f�4 ���w߬�`�E�V{���yyM[��sc¬}�F}�J1j\��h!%稚�����vxR�U���
�u�7��!�N;9�����x+l%dD����1Q��#�(�?�vtj�ky�jKC;!�����ϘlA(�B}�|w١jb���U���/��>�9Z��?b��1�D�=^���W،i��{��f��܀[����"��3��<Y��O<m�&#�OD��8ۮH� "�cr_�].H�^�����,��L�F�D���t���s� bSs[�:gbR��1MhA�_���^J\�M��_A`R���r��:�����%`)�A��X�v��c���W�]�і�{*�����ɢV��7�i��>�g���͇R�z/o_[��\���^��̆����Z&]��#F8z�\
�G�z�9t4�g%����{��P�ֹ�N1�>c�B�(^l�W;�!��j[{7<�Pi�I�z���8�D9+or��0��4�D΅3��ل��V7zz��7f��0x�c|>��a�}���ȣ�Yڏlg�{@�\^}}��ZC����XY3�f�_��-543�}u$S���w�h��,��4B��'ϰ��+�s�{2O0!)9w�5E�~ūt�YF�M��4�,\�|4��#��P	��� � ޞ���~���k�ˀX���3* (��7s�-�|��
	D��c��X�}������W����릘Ԁf�X�e���_>�Iؖ������ �O7;{��i�0f>��G�>�g^m�gL'?��;���5�5�����`�w�o�"�ս���Nr���_�]5l�n����,ĩ��G5L$�x*`��Ӎp��f��ŋ�ho����Eg��j���TF�H�Kw���������o�ޮg�w�?.��'Mn"I�݁i.�)݊b����$���C�K\ <���'xR�Ql�}���g	|@*	:�����E��sn���%Q���;���j�tVG�/��ƷV�R�����~ᑳ}�=���*��'h5~zzLM9��j�����x�(a���3�p��Y������	�o&s��0I��c@
c���U��_ʭ�A�:���n�%G�;x���:t�"q����ͦ�e�c��԰�t�=�|g�G����n�(_���E�<��1�% $q=G?^= "�!Ӌ��}���"8;s�ը4�M��k��|Una'+��Ɂ��O��P<?���/t�6�6>|b���e�jJ��7��C�iFQt���v`v���Vc/���*;���O��iW���P/`�&��(ؤ)ڵv|��(����"~U�;N�\��&c�RpF����<�]������,�ґ�X*�iC�7a�X\�D�KW۱f+����f �`�wl�L���B �/ie"��g�fW�4>)�n�g�����$<0׻eE��[���L�� '��j_Q�W�.�+��lÁ<�P^Ne�j��!g}���F�����d�6X�L-�k�����s�V�9S`Ém�Ք��
���`�=�Gr���m�s9��IQ�+�,�����ݭ�7�E�e�2��!�M%Kc��~��YG�N�>�T��M�M�Uu�j-���/� 6��,&5�@�9 �V#��FV�_O��g��vW�(�)�m	�HUm�-� ~cM�ǿ��@^�G����1s��� Ac�q?%3��x%1��rt��|����8��~��6��Bg4Dmk_i4�V�p��7K��h+�g��<��hU9��U�e���,���E�O`Y�&gw'�y�"���x���dY�+Y6gx��Y�dN���V
�=����{qPI]ڂ���`^��
��|�ʕϛ2jeK��$�/M��XZg����٠��_���{!#��-ԶN5���8P��F)��2�wJ���oM-l��c�~��a���96Ro)�E�i�a��m��k�@%��&4�5bL��ހ�j�mq��&Z�E�&�s������z�D+�{fl��|,�)o�� +pxB3R�A�8ז\������r�;_3&�EXPs�<j�@�t1�kiZ]���|��z����*qyk G9�qo����y#Gj)�KO����r鏉�y�;8��n�@��zn�>]}E�<�"L֊C�n9�k[�D����c�j��TT��7����:1tP���?�s;%^`��}�@�ES�>~�N���v��fܟ��u$s��ň�S�՟��U��`�xaë1y���v 5#s�p2�²�x����Ƹ��y��I��ꙑ�́��dO�w=�:ax{�Wn�[&�����ѫpӂ95XԸB��|'T�bޢ͙J����%���=��T�C:/�RJ-4b���6|Z�~��Q�@�e��u���I��S�E���$�m��ڞ�iۜ����U�jI�� }��#� ��x�T�]�s�c����^��U�}���H�&yGTWR*����ގxޜN7-�PCdWEa1Lƣm�����jtH�U�f��z[ZBP�����Pb��+)��ʻE^}����j9�G�4��A#7���-7N"�7-���@����EC?�h-S���sZ�1�j���Ш+C�$=�.�a��$K����,J�I���u�797S@OI����}9ϒ�N-[���X���1�m�d��n������#,
�}�'�5[N6�$��x����n�ݑܞ�E����-� �O]dڹgO�wˏǩ�ڡ�9�ne��������I5M'��*k5��$���<�h�8�Y���}k��ѐ�4F�Gn>_��vb󵺐SSC�ν��dt�t�a���.���ҟ ���Q�#(d�����5���tA��dM~lO�t!}���r����Wk�U�.N{�U�T9�%��� [���z�Ͽf]�>hв�>�x�i��Q�ok������C��3����.�
���ssXwg<Cw�O��g1x|���N2��k��ޭY/�O�U&�AĔ��)8D����<N���&бq��w�O�=��e�k����ֈ!�w&v��'�o���?��2*�eY���4��wM����%X��www`p��2�08�s޽o��{��Z�������Z��Y}<�U��1O٥����Ɠ-2��:2��(k�d��CF}��Yi�� �p��	�\y��r� #��/��s�O���ۤ��I���.��?4�sG�xy�?Yc�ϓ�u��x6G���,0����ZU��<:1.-�=�r�������_�LJ�#�ć-�j`�\�k�aчK��Ixp����1ܚM���MNP���_e^��u,��W�yH��a��)�ԧq	P�FlVҕp�T���f������:�Ϙ�hӫ��L���$om�����ݒ�?���<.%�v�.��ǒ��',������ߍ��	q�yo���8 T�����'W�wH@��Z�k�͕u_�<�"������>т�b@�ǖ���'7Mb��V���v��삭'Κ�o�4������['��<|p��p�B���J>f�]6�مfߞn���*���7�eJ�p�Nvſ]�fi�?E�oIo��NVHD{���0V���g=@&�����dc�u�%��>�Ԓ�q�����S��͙W�� M��LE6zW'�K��7�����������?�h������%� �����U�"0	N�j��T]���J��0k_v/���y��
�R)EP�_���~����VE����#zׯE�<TjUx��@�=<R4�-ޚ})�Rl �e\��-��X{`�O�d�K7�Z��������
�8��RH�6�ϭ����k������:�x4�CH��z�1Է�(�]	���]��m�5�x�a%���<#	�fy��]�I���?��:�����aƌ�(x32`䐣<c��|GI�4�y�����J�)ls��p�'��'U��'ʂx~�^�<�|q�%hx�n�؟)�=�u2�a���ކ�WC6�f���0x�,nl����z\=7c�R����@��L�ޮ�]��T�t��UD� #\"��篷.3z�`��D�t�B/�pQ_��Eg��=��_�o�>�\�ڧ���G0�Qk|�pO��4�Ի��y��0ko��X�p�~���H�s�'(��Wȓ�z=�ﵰƿ��������/� �^�D��[bN��[oX�с���8���k�ҍ�@�"��? Gۊ3ri�*|���6^Q�� t��9������:�v�t�v�l�~�2�w'�Z5v��D8mI�i�}k����u"��{��7W�a&*����z���Q('�K��㥺*(�����
�#V�Q����/��"E:Ƅ���}��q�L"�5�{����Rd�0_�`��L٩ԑ0oP->�x�t�\Ec����)�)9eK"����H6���pq�n�o�c�����"���,�'��ۯ>�П�d��w�0l&|�0���[��su��z��޵J��Qs��d�8��jO��g7�#q*е�ia�<�K��]/��au��g�-���!�_\d@o}��3oԬ��B�OGygLm8��/ �iZ���9-;�2P\yoW�P�m��
�Ce�6�+�^F�}����Ԧ@�ċhR��G32���L-6�W���~���E:��O�@b2\sA����0�~�~W�N��ش���+���ɛz��}Q%�Ll�Z������&e�H�l���Va���O�������?� ���&��~���c�;ikR�U�;3�؇O�"5>Ay�@���Is��	�"җ�s��:��R�Z���i�ٴ�b�EV+&�'1���D�	q8��h�/j��Kl��9$ɴ_���S�P��{m�#7��ev\
`i/�+]\�������~��7ޘwI�8���W7��"k�m�o�7!� �Չ�TO���.�ÌO�K-�����p���
iV����{$�7�GQ�E�׹�"��t Q�������e#��?N}�t�l��8�4�4�D{U04貨Q���� ���ї'Aa=U��K]T����������-�':o��d���$���#�mbߌ��k�3ضNq`��d��b�j<-���~艇����}ލsn��e�g��]�r�·����d�
ݪou7
`�JUE�h?��s�Ό�m'�~6ۻ[3ɋ`:����<�/��I��%��9F ?�v�԰J��7ɩ
w�KF	�A��X;���Z	�*	�6��X������j)0�7����W7}�����,-9ᙋ}�#S��q��,/��P�[5�X����8{�wІ���ӈ`���3ԏ�3 z��xq7'�>� e;���fOK���hkV<0�U.Ch�f�����Bܞ�WO��� �=��Βr�a:���i�u�%��x��Å�O��՘ZX�>V9Ay��nc�p������<���������O�z���&"����a������$OD�����[�@��佁���.�SaJ���·.�.�qH�ѐ˹�����e�P_ư�36d&���~�[Ԙ��v�ed����"f���B�S��>�Nݘ��~o�w
0J@m�J�*ƌ�%���:���ۆ���0^t.	�Q�~��R����v�j�z�lzr��Ӱ�fϛ�ay�Y��/�IU��-�� 9Z�� :����BP�?�A��8t��{n�߱2В�_^^.�I����˿���P=��n��ZV�����fDU5�in[��(!$d4h���]Q�/�(�9�,���?��&�JQ�Ǎ�)�o�ɚjB����R�kM�Q�u���C�$�}:L��{���B7��Wz��s.�'"�&S�2��Ot���49sC���r?Q�u���D��A謾ؿ�~Ƿ�N��&Q��97Wg�\ <|h�*ϔ0NA�(��1NK.&1������{OB�7e�v
��	j��f��)4��H��g�orђX��P�ZZ:W�,���fw�ԍ_�s�h����rk0�e+|:���R��Ǐ;P�4��ڣ]ĩ��#|��k����=L��}��Q����46�Vrc���w��3�q��#j�V�g���d��|)�3�`=n���%
�Q�� fVʁ[�<�7.=�+��Nv2�v��N\�Co�\�eOcۚ�w�
���'6�_����
	�����J�"�?���u=�d���0����S'��mR.��5k�l}g������ԑ��%˽S�3S�p�.6Gc��C���^�m�^�ن}:�_<�(�<:s��E��X����v䘍~q|�x��bo�AY�$�lG��6��(�YԢa_,H�:R,&Eݻ���k_e��W��}��������֧F��gZ�/�ɳ�9Wb�]�v�
x�"�ȳqX+"e[��Q�h�#�g�*�.G�/sBxf���\SZ���pwJ�SV�uKךFV�u�e�;ty�@��� �;Qu�J��.����A�a�N�2DH5?�d��c\cWlPS��J��ƾDU�+�!*��r�٥��e��WbB�6u��C�M���J�m�鼉�	bė�΄�����1\��\�h]��=�9vr+ۋ�/�����F�.4{^��%I�I��1�A����f��ͮD'�����>x^\s�����Of������ Z���zt��r��E���|c��a�Y-�S&�Q�Ϗ\N���@������tV�͋�:[�̈́b�_��.d�\�Q�S���JN�#�S۱�M�8|�2>i�щ�/���xZZ�x�ɫ��b����c�o���?MuC�0�n@�0��'� 6�c�~6B"s��`��3�FQmn"�ا"�7|7�)�@GAY���t-�n�G��{��W�o�ԕ����b�jpF�+�Ӡ#��s�򛺍���P���CC#5wz������H�������!�W$b�$0��%Щ��b�ӑ �&=�Б2��������h�-�כE&�ɽv�����ɛ�}̳�nx�?�*��gމ�jlG����E�̳�O�<r�%2�,#�� �����k8Ӛ3���"j����ͫ8ļ�8:^����gН
v�p��tlw�nɝ��m��9'�4ٟ���UV�kXC�dl������P�E�O���V�zR�ʗ5T��%!�.�hM)|��d���L�������:�����I�|�Y���7����$@y��g꺧99j>>cZ����F�
����~\Ci$������G-��������i�6ȹ���-k]����k�<s����DPq��6�׉�b��3Qf"Q��݁��5��ԇ�;9�n�#0� wdh�OG�oYI��Y9f{����9cJ��s��I݃�eq�SP��&�wM�b�ـ�?/��^��Uann*5���E���ݕ�Z:�a4����9v'�b�������0�!�0� v��Ե!\4
�9�>�iECV�7L��
��z�Y��$/ɹ�~@]�lB����_��k�?fbS�1.,����DHd�~�T���A���й�n�����B`M��ÓۚO�l���L�>�ji�	����3{
x.ZT�s�֜��K�Ӝ�䅋E���E=�.�	�e�Md<
����'��O��`5Ӯ�[G�&g��&�i��ƾ��6�l�}n�����WvUzO�v3?���:5��UR�̥=)}�$2#�uRl�w����T�k��"���A�+��nX����2Un'M^����]H6A����#��ɭ�anqމ�֗���V6)�=C߉������x�h�V·�� ��8��"_��Q�ű?P���6��|zO,��<ũ:F��$hg16cCo[�.A^�Q� 0���{�D�}'N���9��V�(�tJ���7��Y��<���Bӟc��gr%��g&��P���=��eehnQ�{�bp��P�C5�:�Rb�r�3��}#@Y�(�2~�R�G�HB6<��E?K�M�-F�G�������)Z?�����Ge�`�"�O���|�7��$*h�Q��L,��'�JL�8L��lr��_�'n]lCܷ������e��r:��d���뤻ݨ`��x#��NX�s��1�b��]BC�|uk�G�3�?;��*���s�l�zC�D��)�d��Ⱦ�̔S1>�ϊ���n&r���W�R���޳\�/֝^��g:}���8�A��;5(
^'�^��\好��38�8x�ll�:q#V0�>!N�k�Y�����K+H�nʑTqSEXq�~�^_�-���0��RM8Z��&%u�9�z�
�6ޜO�P��[��_�ȴ]A��~��� {��h'Kf��$�C��'�,=�;Iމ��$�*�\:��pB��)$[�_�M�Im�|�`k2��Y���(��3B��	����x����#��<KҎƳ���H5�>��bعV�/�Q0�"l�V�M��w�q�`a��TE��;̊�	��mœFm�;]�!�m�	+�� 67��[o����S�`{��|Sh�"��#�;�i�ay���LXBW�뺝� Ȁg��cc-gѝ`0�(2�ā��#Yay�f�W�� ��|���-6揨Ζ��x�b*���@'PuaD��Q��^�,�!h��8(�[�Cڼ��}?j��I�?�琢�?e�x��"aʂ���{,���* �.T#o�n*����*(��gw�16��z޿��Q���&��V��!j����J�}Ίd79����qxī��5����S-�ŀ%gO��-m�+Fg+�ȳ��,4�Ch�w7�um�\R�ċX����e��m�=[�����n��6����~EL����_��.�]�˫"�S}�%��-Ʒ�IȜ~�v`���ܜ�~��UHw&��\�PC���n�<�'�3B����s��8��(o���N̔�Ӏ+����g��"=�,-�SX�]�ø�/�r���&q�RLY�b엾�/��	�1�Ir��M�,��3tM}�j��%�f����z;����>j�EΑ��O�R�C�x�f�F5 ?ugb1���(:C(��,u��,1x�% ��52s[��w�v�5y�w�Dm��wT��3��@C{e�w�WR�&�֪�n#Ǭގ�~0��ҋkD���4�M<y��,|���o���Ř���bT�?$�gG�w%�.y��G4��1`�����%s����{4ُ��̜z�N˽�w��#�%٩A�S.խ"Ȝ���!Ƥ�M��Yp,Ĉ�!��D#+�����+8}�j d��F�v_.�������Ay���O0�6���츦�>k`��	3�&�ߦ�~�j�v�M�쨥;e^�"��<v���9���
YPX��!�.�{�hߋ�*w�m��%�N����YM'�=�S�=
t�K�����f��hG���B�!!��AK�JL�d���7@$�4ͷr���� �?��hzqۯ^wq�n7>#����[P�
E�zb���e�̳,D~���9��'�^�ˣ��<�$@���d�S_	��

���E�����)������ �G�_��Fpn�./��ᜯ�x��DzĊ�]k	kV��i��)"%�P)��ia����]N�)��?�lRo���Ol�)=�S���(*�����wwz��8j/�\y��	eA@RKJW�5����+��v�� ��m�����K�z{H��f���T���Y�����������h��$T���B��.�&��;�\,�.�❑7��p����;߮��a?$��̠k&k;��{]��|���!�zD�+�Q*^s��0�փ�X� Fw^VL_�8��Gx���^�p ;~�poTD˟��s���zk�LS���0��4m��$W�Ȭ7�~&2�m8oa�:�\�nӲ�i�?l���6��W�����u�$�q�G��װ<]�Xݤ�)H$'ZZ-*�e���T-�M�)b�a�D�3�D��e�mε$ꯙ+�f(�N0��|�I}��C]��*b���u�u�-����;o�Ӹ�n!U5���ǎ9�F-2�*�T���ʾ�@g!�nFFV�oc��k�M*���4�ʣ�L����OJ�"3���TY<p��Tk���Ҳ��
�ې�W{{��X(�t��.z?�e���º��;�V�ϑA��י�,r_s#����cL��O�
B��4�*j��� 	��Z��r]�ڲ�`p���jW/�J���mLZTv�~�{���4�M�Y��~|�.o�T@ݑ������N_��g�joä�������V@w��| ɍ+��*��䰑ww�������ځ����mC�#��\<�SU5V����;W!m�MfP�b�A�������ww��/��c�v���E��{���s!WW�~17��PKy٫��A��h ����
�Ǟ����T�(�@����h`�~+���9%�g�=�n��|��Ȗ����375�l��'(J;�����D(O���FD���t��	�P����8�^4�fo�k��'�E���{�H�z���'��k�M�ZVj��we[y���_��`P�=��M���̻D�U����TY����c��og��Fѭ��F̐V��དm���p�B�jn�LM{6"�z}!
�*-ȡZ;V%��e��8���:�6�iE��a�C��Di�D���{^�����k�U�\Gz1?Uk�s>�Sf�R������+��ɫ�� ��t��kG�w��$��^ �b5ܞ�)D�u"r��r��yq��y-KWa,�Ov|�'��pۓ1��M�?��w6D�>�Hv#���"�Q�~��@�D/4�:�3�y3���b��Dѧ1hT�95kX�s��A�>YK���=!]T�jʲlZ�M��Ŵ�k� %Q�k����5�&�/��?aڽ~���UA�15����ls���H�ZKǰ�r��Ȭ��D������-|��<�	7G�N��n��a:����/�����d
�q���)x�༮��ų��	�ʑ���"#/��B)��������&���{݃o���������*��?�q����,;���y��:\\"�ǿ2X�7`����>c�8�:�������ngg��cQ^Q�/��l�z|�5"@�4M���Z�߼�]a�N���W鴚�'7�B��!��~����x/Q��Ji�<�A�4r=̏���l�N�Z�ib%n�d��i�S�
�?��G��c��?wt�&@Y9!x��ɻ��<�C�o�m�/��g���������7�C��A+�o��.Ƙ��c��K�ZEL���R���i17b`pOrd�9��
v]�^�4b���ޯ����M&dj�����re���%�]�$�^`�翛�G�?�p	�q��O�+�Pe���߽�\�@ವ�Ȥ@��t��+��چ�*�J�ڄ{��z��c�>�S=w_G�
h��شȒ�����3��st@�ee'��Er���YX�}=��{�/�^��֑��,u{�[�sMFwջ��7$b�ϘY*}^�_��Y:Q�e������[���yb�}v�ʑ��al��.����\�^??���OJ
 &%%�B�Ǹ��-��t_)�����|/���#Z�݉Vp�+iM烆\�P:�ї��E�5`��,��(�ᧄ�Ȟ��{���G"\΅�X��+EE.�ċ� g�<B�^��]��2��ܷ�䡮�[�7%b�y��P����{'>Y]I!gNb��G�h��O�֪3W���~���6����,E9�]�a��wA߽)D=�e��s�ft~]n�����z'i�|3...p]�D9 �!,!%;y��ܷj;�
�m:� 8����ݓ!�f_���&[����g�M`�B��������5�wTTc������s��7:�����X��e�B�##"g���8aX�B��L;���K���1����.��,��������F����ba1rs�������ϣ����R�����/O�q{����FA����#�Bl,=� ��秖z]]�F�{��܏������08,�ʇGq��,c�/Ey9j����5��=D�:���F���;�`>g���ξgcۋ!���O"���h���O=���Z]vQo�uao��@F�!�YK�^�'�Z�f�p�� �i�P��Ǣ�Sr3��P��1:���ϭ�T�[�/����=Y����p��R!��a5�U���4@.%�5��6#�����Eˮ��r�G�`�*dx��[�Ara;�8͇�W�������z�iy���b��o��
>������-�m�d�9S�`����J�y[�fjVA��Lj�R�jZ#z��5�[��?ѿ����/^߬5+K{��r�鬛aYܭK���~����l�<���V�W��kY�B��j�M����jC74c��Z 3�j��&�˽'w*`TL�zb}yy[��v;�����w�h  �x(I�A+&�5(yY��E@�[��]�񡋄��1p��7�eb
W�����b��5�"oWH�qӆ�y���a��WԔ,oo'r�>����?� ��`��t�Mcʕ���¸��X/J���ɐ�"��TV�QY��Xׇ{PeV~�����5"��#G|l��5�_��:����4��91}a�?�AK}+o/�3���c�(��Y�Oӝ��_��=}!�2Įq�*�d$��)	B-Y�+�[����`s��1YEEE�������)pS����i1���Tr���%�2�S�QEr�ԩ��`�wCv���v�e{�� �՗��[%S&n|o`���q����I8N�!��B{�<z{�`{)a��"#��}$i?����5-g�/z4\�(��e0�4U�N������*��<5�r���i��
��j�����7�z_Č����0�����D�:���4F�a+��
M��'anMy�_K��k��.3�b5O�ky��[Ml�}����
�|+�����ʢ��r�K-$�Ê;�=	o�iUlݔ玥"�)^^����Y�i+���SK��Dfj|�aPꌍ�~�����x�˵W�����~t����C��'i��"�6��S���0/&^/��[���2���ߣ]m��%��������'��Uխ����r��
5i�1\� �ƋH#[�nKF��t���_�ݶ~�r�*��|
Dβ	�Ǭk��Z�6Y�%Te{�h�!.آW��̄gv��%b@�X� ����"���
�3k�(��V�;�/z�ȫ�\��65�������3j�x�Q�>������f��y��N�;����ɳ�9��b3� �~� �O�� �pE�����%��c��l�Q�$����qλ1z�K�o^L���R\?�H� ��N�TK��W����>a�j���6����?x2��veLwӬ���mY��\v
�kl�Ro�jO5��[l�$xI~[g��������m����;��X���f�y7ur��ႧV'�1G���Ծp�h94���򔽬n`�Hpa��Ԉ��U�jPO�3��1��RB����b�>r�2��8`��� tx4"��J\��/Ox1l��Ȼ�d�52i��X�Q��)�u��nQ��
� �}������K�j�vg�B�k�t �zyI��R`>o����b5��t|��[�%2��R�����6Й�w�y�M�̅팦IP�1���2�Zo�e{ڲ���i7Ǣ��ti�X�L�~�G��_�b�9].�}B�U����"�Di��y=���F�3i�8�:a�*/.�O6o����ɀxl_��2�'�P�%������Ԫ|S�{�͟�P�#�;Y�zR�:,��mƩ�!���2�GN���3��h�Ň�{�?q�������L[�#�EZ�����å�ж'����}��U��#'>WB����D��Yvj�k�Z��+ۡFv��<�[#����J�y�H�Ɉ�9ؽ�⛕i;k<N7�!`/=أ�1^�!��O(�<t���{�);�v�o<�6i�pZ~���<muiJe%9o���ߣK(#vA ]�}?1�n���ܝ���3� �c�T��e!�$�u4�9�C���)���&dX��s�.�NZhU=2�+�S��Hm��f��9O���;�渷�\������x�`S0�
���Fe�&Yr%��&'�bnR�;s`�	BSI�y�/y�t����*��8��[�>0��]���:-��[�A�W)�?��L��I���B��Ug�(!E2��O;�����S ��*�Wg�t��J�w�K��jT���È���[��~�S�;��Ӽ*� B��o�4����k��w$��9g�28��K��(1�l|�|c�q�{��f��6�[��>C����bTE�4�ɺܴ:�,]�4	ÞC_k��^��9v4���<��=����C���~��/ȉ�Ny�M�(O������Z%�J��vt�#���������u���N(	��s��m^�ƌt@5l2ד@dn`��6�;������M'�}��
Ο�����J�/KJ,mZ�o���}	�lNUN��϶�5��|�v�1�L�!��oO�4���(,���>�A�ڞ�>o�H}�8��v�/�(�5�l�����T~�c���y�UY��!o�w��X��a�7��<�F�,m�.�}�Z5���1�}����CF�I)�w�q���TQ)�XM�^q]%�ZKT�"abfF9:�e��/�-��EW��Cٟ��� �r��ϐ���X�嫭�P;��v�!�~=��Tș��1��t�Ƌ�a�U�����H�Bl+��������~|�EN2H,�Q��WR�o���c�L {�e!7n9�t)�|�7 �i0�}15]TS!��l>�.�OP��RQ�=�G��Q��%ib�����<[^�Z�N�"�C~�[h��T��o�L�����%�R���(��!�qf�%�����m&_��Xl5J�AH3*���/kL���KA�e}v6JgFY��/�d��j�\&��#+��7�y8����,��R��ޠC��.h����%!L����k�;�v�|ɨ�T=��e�<��Q��@�����y<ߠ�8��d}%P"����p߲���B��������zW��m���d}MM){^B~&�T���`W�����\���-7E�;떩c��:�63���G�!�i�h���*��7�S��r2J{��
�꘼e���縋��Nz� >�گ�CV+$�%=�M�VM�O�v�b���8nQ#N4o�q��"A	��ٙ��9���'W��W�v�z�|a��d�НO���|d�z}oÅ/��9���ӛ����5J��1���!�:N��ؽ�����p�L����W������2~�ʗ���sA���?%ƥ�X��ù*Z��1��[�'�9o`��vOT=��<����;޶	6�I�U��9aCY�Ҽ0%����#�MS_�p�(;��N�� ��q� �;���.0������&l��ęK�&T3
^\��Z鋟�9Q�#cX����v��5 4�Z9�Х�����R$ �9��X� U_��Ni ����ǟ_D����kpI�����3_Ό���nn~M�ݝg����O���Wp�[ao���&��6���t��f�2�X�A�_Ai�o��a�O_�$���_6c��3�n0E|5�c֌K��'�R��'ۭ�v�J���`qn� Ӷd\�uF���Ì�Z��ǣ^���e/W�YF���:���6�sף^$P�|���`0&:�7xRȨ�8=��-��Z�2u�Qk�a`w.L� ,y����S�]л5__�@Ɯ����[� ���d;�;?,��֢�|V-@�ޕ���ٸ��5*�u����@��@���3��2�D<�320(�ÿ��8�:��D�@�U�Q�Pf�=�:����_|w�N�_}��X�1���3>i�:;p�[)3NVo31
���BAb&E����5� �vv�9��`�N��5�/�e����t�Yq�jh���>�j�\��;'����[��L8 �7�m�Ĕ�#���T3#�2���	Ma7Q�?�$0�f�E>�u+-8�^�M�b8�vwI^�Ѧ��ݙS�)w;'G��N9~�D��B���A+����<Fq��\$�ӽ�7o����gI�.������=R��-\�vɛp�Վr�Ncy�\]4��y�V��Ƹ�������z�⋰J��D6x��d���w�E�%�lľ�|��J��󕥼@�>h:�M�]Tg�ݜ��|��}�	�r��i�NdP��?eԌ� B+��8�T8>�m��n�)���f;V��[�	Ie E��"!IBi(��_<�����]�J(��:a�CF�,��<EG2J����M5!��4,�V��WɓN�5�ɿ`ƽ�G�x<�3���D����Ζs�~6w��8�3v"�J
=Xx^����������$��8 �r�aA��v������7���պJ�	�o�M7�����n�M�c*�b �8�⥆7�S�zm����1�AT;:0�~�,7��jƧ݈J{ލ�.:���ᢾ�(��u�X3��cB�8�8Aþ<'K]t�X���g�L=�'mL%���I ��w4�A>ܐ�M�����6{�2k=sq,�ޥ�L��Z��n�����3�5֥�ϳ�Rɳ#���ӝEL��$�����#��
>�d��.��7�rV|.�@��i��35�:Q�>vF�W��v�e��<{�<�W�����=�Y#=R���l
b���e��s���	k��ěز��g`����RCSC��T0��\ȡ�$Շ��W��<���@D���)B�)9Ks0W�m����ނ�9�7c���/J�u��q��M~���g~%�!�G4�3+Ӿ�\�,�g#��`]OD��ðd��nJ�^�7>B�Za�U��~jA.�����*�!�t�	@�����B��v�;g��s7.���?���%��u`��q���*`���ȦE�z~�]QaG���Z�#�"��bn�Ɔ�{���:q�x5���h��F��c����%bTg��|�_��f�q���;�b�!6(�ޡ�mU#_H�;��p"UN���a1H��w}�{��NKy��c�E��6I��j9S���L�v�tx�W�7��T Kf��q��#�r��gK�S�� �¡NLNS�՚��}��$]̓�����ofvEIY��̓����Y��Ô���Y�J6wD|<֩��Wgvj*������a߶��쬔�=K.Ѭf�u)�9f��QM��w 6Ę!��!)yd{�f&���T����Q��v�u�Cv��d��c����K���W��1�A9]b��/r"VN�Փ�<+(��W���	�'��x	zz5�%����ngnf�J[[��j�ETբ,W����n�#������
u����w��HQ�N��}�����}��V�+�����H��ihSz����D�oBkb�4� Yf�#V>���UO��F*��;��Dc�ß�����s��d�Ѵ���x�t�����(!'��k��5E��0�X;����i�EP�nz1rno�o�橸Oh�qT�r�����0%%ದS�Ot"�JJFA��{3$�>ؔ��u@U�$��T�������goR�l¡yǐ�h|K�OL�3�x����q�s�� `2�pN����q��S��;15�v����򥾩�X�̫�J��*vs�hT���Y'B��B_�\m��h0#\(�=�I5�N�1�$4�i��]�꩗X��Ze0O�o���a���9�Y:诚Ů�	����P���?"�(C�w�DVե,�Q���3�?�D=Z�}��mV__�f܌��/%����V�t�+�ݝ);���\f���&�����	��x'/R���Y^��(�&��c�L�Em(���S��	ݤ�Ƙ���(��N����ܳ�|�!�c�����e� G������y���M�R@�x��Vw0��b+��̥_�J���P{~q�����ޙI�=��������&*i0��|ɴD�b�M�l�����!Nn�a�Ӄhvy��zYY�9l"��U3j1�~�Io��Q��0��U�8"�@񫞝w�Ze�JE��Z����l�z�q����z�u';[��,��y&�n��lw�j� ����cE>h3~�I/5��0ov-u���{%VKe�xh����>��D��ZU������l���d�������[�>N���]��>d�m�r���&��X^%���Zb�^K��~���4��]�+�F�@ٓ��
�t����*n���o���G�t��]992:y��J�����d��p�å+Q�U��!'N��p< ��%e��M��78������	��e�d3�@96u�J&~���E�,��XF衬��e���4�H�nş(��8���a#CM���ūfO����ØLg'E��g�V�95�cօ��w��]���L:�f-'���%�4�4Ku���+���i��6���M�������_� 2X���ԯ�#�˕��*.R�_w�.Fy=)����x���ټ�<��N�F�Q�	|r��:��V�8��k����!
������;4t��-R4��G�=��NHص�T���\�'����N߶G����I#a�4�M2].����ɍ�^�����V�@�f����"�茌�ۦ��h%ԏ���lМ�jg�ϛ�"1o���5���XŴ4N�[�*Z�r�w"�?f�ϣA������DŌ���[/���/Z�{F�Y��"dM_wst��O��;A�Q�U���3/�L�[����T�V��5y$
L6��V������g�-?��N���@�~A^���oA��
�[�c��ß��T����bȲ��jpp�H����ź�iI�1YG#6�V'>�������R��%҆I������e�͍��-��;$��f(�`�h.K8�Wű9�C�!�N��s��1I�����g�XR�h�#{�-�D.�:�o�RX����Z\P���_蔨�Q �����?Q|q�H٩�$��ݶ~����U����o�%"�&���۱8�PM�%^�&�)�P!�
����g"�l�e�kʖ>q�u�&��k��Y��c�!��,r�0b<A�҈G�}��+���_�����LR���X��:O|���%:w�,j�<�[�̲�։�o����9q_.6�I�������f�ivi�����.B�S!�#�vT�����M�e],���#�fϝ��<[[��45�����i�����W����XR�?�����)�t�_;��.q���l\�����t�~��E;cC��j�r�%�g���I��r���T�nN����Rl��g<|�o11�V��*5�^엦���m$?&���44�x�;�&|)��%\h^
��b���/iə��uk�Cӄ���T��a7�d?[��ڌ�"����T��eɞ+C�x��'w��!�>=1�k��#Q��6"K(iAԆB�%L�������瑯9����UF�b����9�ڃ��:�#����E�Vo�#S�W�_I�?g��|����O&��~��A�u5�٬rw ��k3|�q����j��Dy3JΠ��������悕4x�����*�Հ��~����+㢊��i�A����AR��i�n���Ρ�cH����~�{����'x�������}�>85Y���^�<��4ﺺZ��!��x2t��v������<�ng�E���'iE����q�� ���z�֕� =@�o���:��2~��t��H����|&D��{����\Xm�r�.���1y�>���Q�6���[�%���ˎ[c`&$�G�TC�?ڲ�ح��U;)L��v�vl�^�"��MB�b\'�g\9�Ҿ���	T��ɓE��kZ2�s�r(L�!�;�ks"�h�9�F%�'P'z���P�߷X��m����y�8�d�DJxM���
��I���V�c$�aa8�� P�p��p�<ݕh����s�7�D�_^o�e!GD謹q<�Q?Iy���d|��f}ԊX����q��E��&�D���	AKp���P�$^�~���yI#�X� +-������5�<�LA!�e�#��L��([l�}1�g��(���Z�qf
�|�����O�$B�`s��Y��4-E�Ќ�[>3���[D�F�n�*�"q���4�G��t��
᡾^*R/m��]����9y�0���:&â���"���:>�k��8L\\��w���W�����_+p��{��p��/�[N|ɞ����h���B��'�I�q?�'�řY�ƟxU�9�gD�N��թnl��&}V$��N�NKq�O�fu��%M��@�?M���;ow�x]��4ȁ89�xq�H�mb%�w�w�����ܡ#���_���'�G��p�1���,:�w�
���]�v�w�Đ�o�9N*��adQ�Տ�"ܶ:��h`!|䠴_�~pZ�;)?<���#�Q���(�#�s�M��đ^P�)e�Q���ф2��G��9��abB�8�B'����,��4e]�fy*�C<�{�I�������i6H�����cm_v���.��\�YK��R9���4�ӛo�ؔ���m�:�;�=�S�Ya�R'�Z��uG���3�����OB��^;1�	�t���bS�wI�ٵ�.�߸20&漵��_���4f�m��Zx�;&�W�>���Idn�З��h�冕�#	���26Xk�bk����'L#ή�$܅�PZ`��^�֢v��g��(C�|�ڡ8TC�����i�I�_
��8�2������t��X��)��m��"������a�Jc�%P&��y�O �%e�'�?�H
?�疚8�9n�ru�>����@я�?��j�]�yL��/[K���
�7nZ��z��7J5G�sh�H�J�Xh��%�N���A���Q�l �ܸ��9�~�y'L�M�[>t�]U���ǀ���'�$2t���^�����mQ��H���W���42���m�B�hT�NO�,Z�`�c2
w�D8\����0���5�VN\�����:��>�}1c��E �M�x��a	�@1\&�t��?�w��[��/(�+�������e_�7W[oE}�䑇��|h�o«���y;�/�9Q%о�l�I����oՙs�՚��!���+��h��������ÞbG�9���w�.�� �E�:��.�2n*�e�i��>�q�����,��5G^b�6���&K|��'�Â(C��"�I��-/�w\*Y��⺣������N�U+&9���t��Z=F�3��=/
+:��|7 [��;ú���ʨA��
8�+<����_�%H���CZa�Wݍ2`�N���
�Q͝�)�Jܘ����Su�~3��T�zgup�,Ǚ�:��X�^ΊB�U�f��;)��\�: Bx%{~�a�p�y��<X�J�U^+����u��a-_�9�5)��lf�!>|}e�-�.�'D
�mw�o�:�t��Ve�a�|!-��ih�U��O�l�܃W��iC
k��W�������Ew��YԖ��I�1�������\��h���-r�@d6w���M��Q4t����W�cx�M��rs��f�՗�g���vc�"�܌�c�Gt���?'͕�2=�-�V�{���3\�M��!߅l�:N���LH���50����W���YǳYZ�ݺj��ZXD��D�rޝ\�o�'����a����#���f�!B5�B��������f����+�BȜR�f���7��\\� ܲ�O����%z���	��i�o}��p誙��9����:T�Z}n9f�;.�&��➡��=�����tr�I�,�t�i6\Ҏ-F�]P&��QJ��o~��6�x8iI} �k��������(}Z�q�\ٿ��QOrsؐ�G:^
>BҰ���θ{$�s1����5vq�=M�L��&(xr�9|���ju�yo�N hѫ�jد(��R� ��P`=68���Uh�a?h�g�~z�Q��2,s�I[zs,^��l�s���2�d0��g�Kjfs�p"���~���(�~/Ї^�W�[E��*����$;�������?��O��L���2qS�`M`qt���c���,�s��"}K�_��+�9MPr����,�q�ۋ�M�e�${t���6?�?�!R�v��I1�K�{�W*����d��z=}Vt��N3(1"Kd����q\��-��H�y�x)������$��T���Yr��l]>���yWm ��i���8Q��n���G�h�1�H�9�XS�Lp�mt����xx��M����)��v���x(B�%jSg�ü�M{��\z�z�5�ޠ(Cjmn��o���m^S��b�x�W�P��q������hl�pg�g%��V���b"�\�V���2Ky���æ�\�����}����#���=i� �S��P��!p�����zU�gp؁�K���w�P�p8�΍#kL�{ꂀ��孝Hroy��i�Q3��]�(�
�\y����'mi�Y`נ�ܑG��}rq���G��:�Q$x�ʉ)d���b}���Wϒc��o��SK��W�њ��p��v��_�Zd�������E��h�8��H;���{c̗���f%���5�Uq?igq���#gX}
���h:�?�:r_OdBŝ"�����;n�Â�F��*ͯ}Ԓ�o��k4�9I\g^+i�����w	��`��gŜ�2c�Y��Gv��1��_� �>���+�0���|Ru��=�>������iʭ�)юp�]����͏\�Y &���ԓy�$"Ku�k��V$����O�x���!���eo}wa.(�3�$.�+͝���^�C +���?�&�J�m���"�{�y^��æ}��f�Ұ $om,��u�Noy�o�{K{Kp��P������9���v�Q� ���]�90"�ӊ�D
����g��4�PH߾�/�wW��|+��>�д%�qJoYZ l����H�:m!�$�@M�5F�����s�i5u�0�A�w�'��R�,��:�^�Y_\�Oٜ�Z��K��%�W��Y����erG������N�?�M,I02��Oč::Q�i~�l��k�Ku�M�g)��ﶟ��x;�A��n2q�$�`S!M#���}w�z��b��gH���?B�Ѭ�e@ۖ���������\�Q{�|󾰦�tȐ��(Τŝ4�9�#���g}��H��R�w5�����'pĳG$ɚL�\g(��O� ��5�����m)��oo ���=��K/u�b�VkL��W�ݨ(�Ѭ0��_�Y�م�ʘ�W�*0dK�)HNU�R��6����Y:���#� �T�����ZxVU��{E���rW�|mP	�����6��x�O�T�����Wp�n��_ `���&�80�=�@����d�,�q���X�o�,��cdd,/�n��V�uy�t?4<��o�l��[�N��*�ON*,#o@��s���IGF"����'��*�Z)��
��XF�p�Qæ��e�8����[�Q�����q����e���jF;7~3wq��M-����]Q��Z�˄�-�~Ԏ��n�e�R	֨s�g�^��BK���TO��t�l>���
:pワfJa��t���O.�:���4�.~��7�O�(�= 끝a�O���w�kG7q�E�ͫ��;ӟj��/x��J�g��v�+LPh��.G2Ѿ�A1_zN��������d���=a?���Zjb�����+#�v ���ld���h��=p
��ʼ`��a�\Z��sz�����yu/�"�>E�y�-:��h�54�Il/x�J�;/�y�uh�|����+��5]�37?#.Z死N���(���_5�g_�ϓG��?'N\6x]��5��u��sd���	�q�[�r��5���g>��F�u�08�v�� �̇5��5�i���7�pÄ Lqf�h|��C�w�"�Ln��-������)�:�h�Ȉa~L/��ƬgA�)�y��,������ǋ�� �j�&�y 5����&�ro��'�0a�/"Ɯ�z�*a���8n��jJ�iK�hrSO�����"յ3�%Na3��=��[���8B�=����P���v������Xp�[R�5A�cε>As�`���4C,�3���yߗ��Fy�|��� yZ��n��÷c���U��c�h���νG.��O���ˣ��9�6p�;��������{��T�å�a],L������K�_�ž�sQ��x�
�+����������sX�V_{�F�J�%�R�8;����{����V�ǲ�h֜]]�o�+��s�$�ΥI|�[�ɔ �nb:�$T����8����E:����/|<�﷤O��F�<��{�h�	�e��&'(�	e�z4��a˫:�x4��2})F���Ӿ�uM}�9�#^NZ�C�#��q0D�ʛ�����R��|��?�fi�w���bi�պ�J	���2��rH��R�Y�"ȂC�<����f��F�3�3d���0D�ʏ:�l�����(�j�̚w�������Zr�Ւ�4�s"�;T��t�ȁ�¢��s��:��]�a1e4��v������{�����2�r�e��:$贿(��������ܰ��p~<�[���i��Ag_�;����(��%<�Bߕ��'Il�L1� �D�ǐW��J��8�9w�'�_�{��c��ۡd'8���l�o-(<����+ �ƴ�����\]�=�G��A6Գ�!��C+nt�J�\7(^"�!��B�ʣ�bc���/Bt�j�s�vs%CHY٨0Hy������;!0����DCC�ԬG����("dp�$�3A^�R(� UJy�nW<so�.�Д��,���Ԏg��L�o����×��U�L�߭

�����RT�*x��x~��]���W��B��ԋZ�/p.8��'�2'�߬����-K�J"x"pj6�	ty��E�V)р!ӕ&�ګ����C��v)s�;��?1��W࡯��ƍs���scaB��"W���ǆ�u�n3� �!�ki��{�z�>�jI6p�5�@��N�_����Y�}RO����q�ev��(X����~Vpfn[�oE��]{Hs��W���\��+�R��,%w�5�z��C��F��mM0���Y�A_�L�ALk�B�B:����KsV*��q�۠ɾ��'A��n��#FU�mSO�F"��v�����}�l�EБ�}A�M3�,��ID�˹�n�[s�,�
Ϟt�����+��Y7�bc�Tϱ�:����/k@{���G8U7%}_���9�X0��n+��{�Z.L��	%��M][�<c�&^A ķg^�J�C��
l����x��*l�����N�b8��r���UE,#!O1)���[u����m����]��"��!IG�_W�+�A�ޅ��+�����T.��h�7��	�4�{J���8����Q!z�z��>5���2�3�_;��f��,��L�{ɬ�K�@�_݋��7���ɫ>�u2��ѵ�om�z����A��Q�2-��7ڪ�D%J���Ԁ0�/Ԫ�H����'Y7�w�M�Lף"��'�E�Z���)��M��*lW��h�H��n�����4�&��Ξ��aT��Ǽ�s��Τ�q����B
�']�F\=�J�es[��yM!�����hD��x[�K����[R��O�b��E��������]=�t�G��j�S�	��;�	���"qzz��`mpL?�r�Z���D�Z��=}�5�nXw�2ex��J�U$f��}}�n��Y��v��}L��������U�<'Սe'P��������P����ٸ~�̷H"Φ���e#.n�Br2͂L���t΁�a g��[l�Q��g򙮳�(����Z��c}0�;���x��6��}�3����v{p~�*	���	>xVJ���cW��\Kj8%O+����đ����0εpi�V|��נ$����7�KE�Ώ��]KY`�b�-u�8�4C���RE@&D`AM��S�p�agh�Wa�
z`�E�ɷ	 ��́�a�h��\��z{�b9��ܫdޗ2��\�7
h/�{ng	_�oL�C��yf(.�0Kʙ^����m���|aY��0�;t��ǫ��{���,�;���n�9��
n��'\,�[Տ��4(��:�)4{������=t�M��B%
~�՗���|\=�\*5J됈��.5���H��L��Mv��
�j�j׆�:t4I��?�����7��	r����9�"���U�������2CBP��$ߓl�ެF���#��fz|!}|���[���2���?kKP��K^׻
���y��ez�`Q��un~�ޅ?D7o�dԨ�h�"|��b�w�u%M~���U���Z�J��4�;eK�d�#�\Q�2�b��ႁ���X���FȆ���,�����1:#�����+�=q�4x��/\�Odv꥿'gm5�c�\+��W�{�9S@`�0j�9�Xf�� ��'�ieGތ������[Ys>'`psm��X��.]��lʖ��唝St2�/?��ũ 3݁�[�wpk�ܖ���O���W�w2�ó�m��U�4��9)?%�����:� s�puL.���ǽ��&��H�6Me���������z�g�	�lΊ��Gq�Xƿ4t��C��*|XI�2���1Y�;�]� ��"c��f�k����'_�S���ܖi9�g��z��f��8V�M��Bw����>:�Y�a!]ܭI$����Q����a|�װ���9���[
���U+���ť�9�)��xH��TX��!�Z_c�ƾ�����'��tڿ��e,F�?���Ei�^X{����Y�P4=�����Ж��,+�c.���l��/�g�z���.H���"T����/WHj����W)B���L^� ^����ꔀ1�Q�
�CH1i��O�/I#�r�;��u��+۴���1c�1�I�R�������pa�Jٓ2f�#-��#�V�'�_ X����-,���,U�{D�v�l�}��(+.�3����ݗ�ž����Lq�Ish~֚K��H���v}�Oy�cY�/Ԗfй"����6;+bC�[��_3{�I��g�V�$u��Q�+).���+��I�KA���p����s���g+�]q�?/ �"��3��������W����d�??f���s)���^�� �^����I�2y����7}l���A�)����Lt�z�ϛ���EEÝ�'av	~E�4��,`^N����k��D ��ldB/岲����teW&N���p��b�N���Z1C#&���l(��~�ܱ
��#9�G�z/���220��B%��Ľ�޺o�C��-�W��C`Oy�/�9Y>]��E�����L�[K{͚��(¤ˊM��!�_���H��G�m �-�+Ya�$2���@:qgU���U��(�i����e"�0���͹B?_�6�J�d�?=�\7&݌{1���8m5E>gҴE���,Q>@� ~�(��K�v��:3ʭ>5���	i�>��3x!�OR �b#~ca��6�e®����_�fByWH�M`C��`�u����᷽{�y�0��{��B{e�s��GS�6/�4#�"�U%�]��;]_��m(���>�˒�0[�A�O�R�K��˙�"C5�;�ݭ��H�b�,$��k�dɸ�ￔW�!%�0��i������s�v8#n;׬9������O��z�uT�(�ka�y(��1��ń�lD��|jr��hn�OL��w�B�N�^�ь�A���uIpr�ibQ�p6b��� ��E��E�SG\��BºT/h>ǥ�o��b���y�Q�w�q+��!�����Z����P�t�G@�v�Q])��*P������ޥ(k�\@��+�;�Q���>�GQ>ԩIG嬆
����1�LT��6�[(��͗�!��ƺ���B�q�>%p�����.|�� �r��=P�]���s�_,��sp*�I�4*��j��l0���z��"�	��y��Ys��;\m^?ww�]��>3r��&-]�d���G�8��u� ����q���_�Ug9�i����������ӿ��C�_0~ëL���}����J�l���$��&'t�`j�/�~+�ޠx�	f�[�v<��a`����	�q�`kҏzE�K4ԁ��/��!����H�f���B�>��W/ä�,�
�Wї�+|��B�M忘Z��IĢt����!S����-G�/�˲��i�Ҷ�n�T`)��ѮWb�V��]���P���9V]�<F����7�j$�12~��v���rm��{�����
	v�E�K��D����I����bLzGm�tq]:����^l2����BC7ʹj+�R�������z�J9�!�L��Ce��C����l_,*Sm���h�]�2a�cũeM6,x>6��o23����M�n:^�vj4ۏx-��!a���*;+�����~�������1���}7�1��.	�GIKƪ����N��O�4'�(O"���E�û`��w�j�������v�p#��+FNt�֗��5g#�@�LϽ�G�h]�� ����:�� ���F��K*	��s��P;禉�Zd�(���¦z"��8��P�����m.�>�����ӗ|uwf�h��FCm�K��}��Y�j��-�^#���E�(l^���˃�e^h�[��Om�:�r<:�ֳ�ת�`a��J�}~6Y!��s�e����>���8%Ӏ��
�L���x��錒�5�GJؕc��o3G�o�D&F����K������#V"��߼l����}�%k���4N��HsVߙ	����f<������=����9�B+��T�o�*���d���(!�Jw�\�(8/�����N�K�:J�LT|������&�T#m�`����3��߈�o� κ�,����|A�]�_ ;w�IdP$g7`�͑����:3�z߲�����w��|8���!S�� ������g���t�Э��vd�c:�Ü�<��|8�1��+1�������?�/��V�^`y�l�'_K�?�p�W}�B\?�гE	8��|C見�����_"s'/�.�D&	����m��䙺����(��nU��Sa�9�JZC)�Wr��;���*z���)X~oQ�4rư-	x�p,C����!vH�E��]a�6�~�����oF7|�Y�i�%��TD�BZ$ɷ=|hjk�Ƭ��+J6*V����ۦ�Am(����F����?�^�>:�mSD�hR�v$_~�!�
�͵9�u�L�L���!��;�T�JF�3Ͷޭ�dk8>����䥾�՟��p1`�_�z��]ô������.�Mvhh���+.��׶,��Ԥ:a�
\��
h��B�x��Y�P^�UKFp8�����lT���0���ǈ��O7��a�B�ث1_`�� (W�������fK,��g6��w���ërj@��a�_5Qb��<` ��;��B�
�+'3������O����w-Ch��׷��|��.���������b��S΍J\��.4~nf�<��Vn*e#��S��[�ܔ�ϫU�/C�}��Y�@T������3�j	4
�T��cKϥ���Ռ��G��!��J�P5��� =W׮������/�u�}#�88=cZ�?k0,<Gޱ�}������='����<�ǁR�zwk�M�c�\�
q�Y���6#q���5ip���.�vY�/���םYy�C��:�YT>D#w�#�r���t��"��������wBW��*VG��b���<%�GrH	C+�1��՝�j�����-�"��;�\�c���WHi����TL�����o^0�#@��K� �]�ӑ�`O% �S�����v=���R^̅�v�-ZK���`��H��\�>�vl�:n���G~�z�g0�3��=u=j�Q�n���e���>���u�q����������診��7�xc1� ��f��ӅO/oMm��\�� ��Ŧ���=Z�S�2�֧�t[�D���yZy����Α����8���O$jM!5 y��5/خ5y�1�x���˓�u3wp|/%�2��8�r�᱉�V'����?W�;n&;Y�W����E���:s'e$��"ڲ9���7���yeI)�������r+�(�P��0���5�	��Pu�#���N��
"�=��t��~�_,�ͧ�Z�UOX�P:�����m�Q�]3O=d�]���?����+F�d���*Ā_(�sz�����c�м�S
I��b���O��b<�?uy+|,3����?R�=��K�W��1`�oډ;��=�b��k"h~��{����.����}��NGJ�s7^���3;EpKJ�V��?�v_Sˌ�l�G��,�#������R��H�@��+3��h=}$<���'��4��p'a-���I�` g�#���Ou����f�g=@�R��.U�z�W�U�]f��G\�L��X��������X����~'ag��@h<G߈���XvӲ�i���4�|�j
Au������v�k~�᥮e���0o���Č]Uվ�vE_}��"C��d~ZĈ�ľ,�a�E��~���3�����hN���K����f��p.cv㣤$����<Iέ�/����{�}��|�<a�!��zR-�d���5�*Ns����v�^�Fh�<�ѿ�<ǈ�8R|��}"�����I�v���Ѻ�	>�r��z��w�g��e��@Eпu�����~dg�y�,�3b�~${��m��u��Ni|xɿp4��I�O�?� �<ֹ����#w�fWLv���/�S�|jJ���@1�������p�o�o;|q��z��d��yy�����f�(�7�^n���x��v)��
�)��?��Zoηѐ���=��E4O������ܵ"�\i,�/��|��e����"]�0~Q�g���԰����suo��zu$3����{PaT��(p'��p��w�0_ѫI����M��F�VQ�Vʞ��Q����m����Ԅ������t�����8�=�����5~w��anQ�N>�3�9�,��6��HA�[k�����+���������?�\�A����iȩB��O@�5wl�k�Ș>�]��߽�kn���k��D�#�������w�N^�6{z�?����F
�~j�;��bm�oaz��N0k�'�@�v�L�n���i9�FF���l*_���c��r'��_p0	�J��N�{�S��ȕ�8�3�w$�k"eX/���CU�������+����*ر��Y���X�g29�-�(`���]�]U7�;���"�y��	� C��g�/��(B��WW'E�\��m��ͨ���� Sy�6{�����\����'���q~�3#٢0r���u�/�s�c�������b^��&����ĵ o�֋A~`N�٭;��[��������fmR���+�&�;-ڝ�%6�+�N%�xw��|���>�ݱ�PZ�>����\��}�6%��ȳ	�j�]� Oqjӱ����E����ei�ØK�t�:6km���C�	�i=W���Ur��A�^a���"6xZ[�H]��I=[�<,Vʜ�$̬]i���eK?OWr:����A�J��R3�_���~v���J~�0�z�����f�\p�ɹ*�8�^�'E�N#D���W�&ƅ�%��]D}��i9`ڏ�W��q���v\� �1^b�6�/�t+����S��q+��\T֐K�R<�NGod�����v~C���|P	.I
��������=ۙ}U��B�K,:���Gұ2�W�M���Ib��>�HX��h�F�W ����K%��O�4w`4�������n̜3�r�(���wF��Ե*m�d�h�홊Q�N�${ؙ?��c˻����/J��3�7�7��:~�q��������qH;r�1T(�9�qC��kӕ�L�O�U���$���1�ӟ߆\�����؃22A+��PU}��L�_q���/	�BNs;�f�
�����|4>⽈�@� (<0�g�Y���h�V�Vb�}2r+J����сy��v�k�\vO�N@�W4;�'#�,V���F�ƞ��s�A�o}���O{	J�2�#�K�_���H+�� c��[C�I>̨MU�pX/��[�h�8h�/o�$�K�GkfȢb�5�ufp��6��9I^-�~��b�D�>E�ͨ���z�u�LM�7U�}��Y{���xap>��F�����)���XU�q�7��7
�A	��6j����It��5�}����C�����e'd��Y�����Ą�JB���~O|n�+O�/G�ca4	Hu/��S�(}	��#�ZZ���u,�`����Epa`aɧˡTL���}C����48�7����rmF'�L��c��?[>���u�:.*Y,��:���0SJ�˲Li�U�3�ඈ���lCy7�E�Q��F9�c �8�@Y����G�꿈�@���'�-��J,{.��ݟ=x=�C���*���$��[~����G�T�}������#Qr���^;��5�~yڷ].��WV��_��V"q�8xB�	0�؃w�_g_�8i�d��:~�Ѕ=��&@�������g~��کJ�o}�$9[��kf��2,ϸ���|IE�egΫ����\"�T������J�T(b͝,���ی��\<��ו#\�)����#cy!�Pz�������__��~+Lh!P��i��Z.&��E�+5h��W��c��Yq#x��#�x�%����n����μ��՞5L�|�k�O{$KV�	�T�O�0z�	�}�[�U����(}_o��U	16���xyt�2��'�m�I�ʡ���=~������2�7���B���X�~N`���T���������1���`�$ �l��2!	& �����:�MwlC����%xo�G�rGi��wb;�1��(-���5Q�7u���~VF�o*BX
JV'��o�ND>̻:��T{H�ӻ�e� �=�G���N�Ҿ��H����ݘ���������p�
�t)Q9͢;y>����ނ�꽧�-"�9��o�5n��:F9�A���o9��d^��T���[J�J��dINVBDx�W8�~\M������j�~Y�������=���L�?�Kz0�����d��NN�&7�ݙ[� �b�L�K��\�ZL��6��F��y'u~�s�n�� "��U���c�!��*�N�:;g*:[[�`-�T¬$��)R�T�y����PO,�T
�"x[ZwKZk$�"$@��	���8SVh�����.5�\�]��5X׶�>����|�^�R[{}�,��-�!O~:91�Wۇ]��m��m99��67�r�?��o`[���d�̻g�7�5��pk����:y�J�� KP��ϓ�IlR�u��?���k��G���g1�8�G�i��>a�牦���H��V��2�d��G:RP�j~"����vm�Ej2u�k��&4:Y������>v���9w_�R;9V��YQƸr;�[�+��FԀ���Z��Д��^ދ-��%�IrH�e������o��16Z%o,��S'��Y��tߔT]}UC��	��a�"�^6���o�q�r�]7�����q����������*M�i��Ǵ��#y!h��^�"hEm�VV�!�w���t�>�<��b`VU�����~G�#��&ݳ��HT�yI>I$�E��wPPՂ���qI�2�bH����kK)����dco^���}���	�.�d?qX������|�a�
��B��`�2u��|w��cގ��`c8Ѭ/�<~��ݝS��҄����M>�m���U���b�e�e
��
�w^Г�8~�_�d�)���o;�,�x�p��O�^d'j�^Fp#�8�}�CD,B�3�XH
���hB<Z�or�Ո0<�s���G�e���`忪��F�Ye|��*>��	ŔVv�U��N~��&�ӊ��.�l���{xd8uh��+Q����*-;}�ށ`\b��r��74;ƚ-4�\Z+��݌���� ;?�e��n a1�8�d�/�pءU���4�u����sYef����J��$վVpx�+����i��
�g�/��_���80���ʒ�1�7��y1�
{A*�`�����N}���<�7d��e8d��y�3���9󦼲�{�ht]���(>&hOc&���)�M/�A�e�6yِY5?U�N�o(��Y�?qE����z�^Zd�9r;r���Ԙ�g:ä�%%-y�E���>#��)����0z�$'w��C�w��O�f� �p�_�BG	{[!��^���IŶ+�g���یo��>$���N�=�~*c�{�&��3�sEN�m�r:n�U�(ק/��u��Z�;�pt�LU�`*�WH����7��l��٦���B1/��_�1h7�'�������^ǟ��>a��sn���U��\�<	��13�4ӫH!7����FY��(N5[���.��8h�F�?Y�����̪u��*{������3%5zaNe%����RB*q��Px�wt�>[��9���,+���ƐӐG�фP����MT +���ZGdgy���N�?����kN~�CMU����D�F�2�Z���R�|}��i?�k�7�P�PX1 �2���,��@$��Z�m�{;�ӓԸ�G�6�K�-��hW�B�Yk�̮��>W؏�$��q6e��Z�zZ�(����e؁OfN� kY����$��mө��I�a����	����.����KoNT��Ex������a��\_����53� X�ڊ���eI�i71��xb8�I'+���Pu#@������z��s��w����}U㊇�N��O��|��݃�c1�<��zH�l"�w����/�-8�
�t����yo?e@���+;���h��ɳ;�ݵ�y� �UwY}vQ'꧆9�;Yd��1>��q����Lrٗh5�s�$Z��~6�~��a���5��(0I�U�WKF)�m��^�!�Q���۝�	��R��Ru��W�p�ѼؔhF���5�t�E^.��䨺O���l�� �0�ֆamEy�F�����)׊����ţ���J�/���]A��+(���Ifא�}~$�WA����Aб�D/�L-404Tr�bE����n)��aR��d�P���Ô܅ն	���cT%W��$��ɨC�گ�������e��pŻ���G�����p̲�*�R]�ɏw�8--�- �]�(�����vR I*��-��۶�����_˟�/�F��7Ӊ��*�b��ЫM��[�n�LQ���e�O�]HP`l�#k��=��!"�њE�Vc��[��
z����A�ݖ���7Lpz�Y���T��;���N���h�@�:��r����7X��Ũ5�w���N�T���>��05�#�"�'J/5�� ,�}6+��de�S�hx؇���LA�x�1�#N�}%��8�T"��RHց$� �N���6���AtHǛa��;jy%���q�-ef�������x�dK����1��z���yuϳ����#)QJ�H��$9�n�r��w����p��J/�������l��C!4[���������"����E��I���"r��rP�q�G^4�h�/a!*����}�]����^�g���F1���{Yh�1ŵJIRǢ��~rp)?謚��%��m����S�ō\��V-�[��׻s�/��P�
B���1�����^���^����|F�~�#[�ڮX��%��/}�o:�15���B�Fe�����	����;��-��\\�\���w���5@�qЉ�4E�&��2=!i'�7�}���PFpY�-�S���[ed��3*{:���=�ȃ���bSȅm�*~s�1���!S�ɗ���܌����oՙ���.Y��
K�D��;���Hp^U��W,�`�|�2sс�E�O�?D�b6�kXT��\UFN��8�ճ�t��:g�Xd��!p���#� `��Whq�잫A�l��7V�\$'���~�S����)P&���\S]T�	e�©;����c��v69Wp�+�u�ܻ�ns�:>a���S��uyd��?��;��{%:AD�D���{����{!D����� �Du��3�(�+���w�}���<s��k��Z�^�>R����_��i7�X��b�� ̗����oлKB�Cz�_R�0'��d��|�Һ�ű�Kbf����d��ycR�5�����(KC]���ᨃ;o}V���9�'�ɯ;�ئH�	h$oe�Pu�H�	qH,��@Ӄ��w)8`������j7
�W��F��r
N���e�����i�KI�+�BLPvn�h��6w,⠗I�?v���o{b�6j�h?�"�$w��Ν�/���A�%���G��ܐ`� S��Z�y��Y,�]FZ	�a���hLa��̤_�/����Y6�e�O�M�V����j$Ҝ����!w�k���g��O�|&����/{D������{��|,�k��h�ڮ���\�@VB��l <�К�i�>Fkc;�z�OؙC�{ҁ��nWs,�����_������,�xĚ�u�ѷR��MZ��/T$`00���68гX��&e��T�������M����CF�gGD��U,}_����'���pUl8��ƛa�9m�D99��� ��R��n ��7��ˍ�K�R�(+�0�t.)uQ�J��A�j�=�G��"~�s��)W{�*�{�L����]
:�#�P]	�O�����{�y(�$Y>�=���#�	ڔ�Z��I�"������;�>.�2!*��S���D��\������t�������D�����b�5s��4R��8jErk��F?oFa�KA����^X��/cy^٬��8Ń�� �Qňͮ�˟�&s�̃T�f�)-����U�[7Oȓ���6������Z�ƽUE�6�z�.D�'�Ӡ"*�P|w�g~�[j3>1��*_�{���z|⭺�y�u�|����[7Cz������g���r�?��
�=V1��f0乑����w���1<�ʨ%�f�O��T���Y��S?6ѿ7Y\�@��ic�;��������ZW��r���W�!�g�s3�z�V؂�t�x��7F���ĈԞ�Ę�Y�o�:��
7���u �����x�5�[QL8j�@ān���Q����%�c�gs�zScq"W��{��K;��}=����+��ܷc�@^��<؃�/��qIe*+�{�y�n��@��H1fc%���1#w$�l!6j)�]e�M��e�a �����4�d���˕���o��GL��,���1���O���8�S/���G1�84��sY� ������٭톺�<�K�R�%�,ύ�C�I0H�JyL[����r�}�]����p�B�J7�KoX�?��f�}&ǵ�����r��|ȗ�R����׫���z�L��P01(���ؿ��~��8@NCe�"�#cr��J�.�%F���_��ۘJ��`�UL���8}I���'��G2ۏW��%�%���#�o����|DÈ.:j��'�[Z�Y��G�D���M��jU�!�}.0q֪����"��M���"a��w��ק�0z-�}�'2�y�C���Y,�?��;��p!-��u*�1�!)���ڦY����I��d6Y�(��^s�{.g !��^VU�.Z������C��G"��7��r�8T�4�ڶ��߬��������j��qS}ı�x�ӋNz�3lk�h�P*8�)&��^^��?�!����[���¼�K��%%��!���%�P� ��&l_���M�m^&�k�<"�bE|�lҿ,���t�@�$�M��I;�����;��q6�z�]-9��*�V����~��aWg\�ol!�ɒ��}��x/��Q��Q~�/��~�+�]�}��$�_�upU��P�Y��&��|�l]�������dK�Q���h|t��_6��Ll��:b2��;�JI56k�c���Y|g�(�z4���E��N<��p���� ��y<���xV���9�`d�3�`DTU�aq�\��s�����g.��I}��3�\�zr}��o�X�>%(�&�̨2���nK��/w٫[����߶<wuv_��z$�4��%�G�r>�OK���Ā"��\|���HN����m<k_?� �ݺ�,3�_��Ȼ�6�������{���BH��D���)�u
7s3(�W��������7����i&��|!�����S�(���اmV;=�'D0x�����E?��ce�����e�c����C�\���uBv���*^��;vn	K���E.����U�>��]�VBC��2��뭶���6��f�����r'w�4-�����&.c���I
��c4���y%��@PI��@'A��|��D4�29C>?5~����L����G�C����AMЙ�^�=�I(s�o�,��p�q��"tcv_�TH���O�9ǿ�D�u&&J�o$}C����^�g�:|�b��<���R�^�QV6�R�4Vu���fJ�'�)�Ljl������O
Q���?���d��g�(}N9&
Ҥ���^�T��U�g|�m�8��𜡆�C*3����"�7}!=>W;Reb��J��o���Du�K���
��P���)&͆>H��k�Z�c�z�$7����C��<��pI�TD���wͫ��������$�L��drBR!���Z�Ĵ%��y�q��(�Q6���u|��l��h��d���~��.D���'��)k��	�^|�����1�.����xUrM���Бez����ْ!j�_^��<�w%�@\�<1F�z���󉑃�5�e�,U��&����,�:��q�0k���m�g$�~Ƒ�%��N��e���54�����s[C�xi��_���TX���|ʓ�0�\�rK�/�#�G
��������@e����1���/�	g��� �V����h;��
J+mxY�n��-�/�6c2��Bm^�!g�[���a����p�'����.=Y��G�^ �J8c��j���􉫇���j����5pX��A��V��{콈������� ��[^;��ܦ}�m=��ұ�P������:�+#��t\˗p���s�."����>m}���}g�J׼����[���ʪ��ߋ���dn�e'N�3���F����:�S��x,/�_�6��Y�b���Σ��Aco�F/Y�*e{����\t��g�N�2�Oܱ/���x�:=W���e-��=�w�~�a�����l�:j,�ok����~��)s��52�H�������ʲ�!��e���(�<�]Q����" }A:TV�[ޏ�by��\ma�� L'7�?���u�L�����P4C��I�H����^.S�s"R"G7�|�G̣��Ot1�eM��0��H߹�'1�RBt�1��qJX�I��ɲR�����#[%a��V��O8Z/�>�� H�󊴼��;�=����YX�%����o�5�t^��m!���i���V1��w�P�y���1Z�֍N���ܚ���^?�pw�����L��]mW�Ww�|O�5�iQ4J�[Y���Y��A,�����X�EˁC�ݓo=m��f�'��q�i��ɝ�ݪIOKN�ڥ.QXgH�o�W�23L�D����c�S��<'�b�wi	�����\sGM�d�T�On�H ��?~�R�uE^�|9n VPN���F�_��Qo-�Q�S���\c�� dÛ�GͮK�ۤ.lί�q?a"�1���b6�\��)_�C�9�zİ���v/��K�2�K�Ďv;������aI(y|���SҪ�jl�7��C���Wi0ޏ���wi|�����Bq���M��⒵�x�ǈSϳnE��R�ՍĨ�.�D���$�}|�&��p�Fv�rTܻ��X2�J�~����D���!����Y��Z�*U��XÞ���列̸[Ꭱ���ڨ�{�I#%����m����@��&K4�������v:y#��Pм.o@,NJU���[M�m�+���:��;��������%Ѯ�o�-�������dc*���NR�
, u��GX�c��#�Y���зҺUs�OF�$����]��x"D}Ե���_��1����bW�p�{"팿U�
�eK���2�J���8$���}�f�����|���+-O����8�����AN�%�|W�n���ߥ+��^�+������ۆ����3/ߡ��Z����[}����4��{�1{n����4T�H�>�h�uqS���@�;��E*�������Qt͊c�q߉T"�o}���o ����Ft�q�k���۝�]��w��\�����+�-W��sB[�W�.��Ydsi����}v�d�&���n-�!�a=ξz���4�����_�#��K�&k9^�=-����7�J��&员Z�C�Wjַx.����v�K�`H	���΅�'�Oեh�ʄ><}'��#���I���ōd�<g�Ψ-,�$į�m��q��7��J)��Z�E�v�q+�����Sg7�a6<��h��R��������镱��aє��l^����M��Τ��e{���Q���bJ�e�@+�����sIO	I6�ƨ�=Ԋ����_�Laaa�G�#��mddy��J��/T�!s@��.zp�!jp���;��mSe�����0�$r�%#��,k=Y�o��-�/��<Iv�Œ�R�Y��Zqi�G��v���$����ch ���rޮ\3��'ui~�ُ
"�,{���*��E�m�Uu4	b̀��v�ֆ�G�-��;[�r]��U8i}����m �d�'ស��޸ܣ�e]w��'�x�;'H]f4��r�N����=�q�r��5���8$G���WE�?!b�,T2�+��-�0|\F{Er֕I[2���)Q�Ȋ�ZB �n@Y�2��K>���,9���dW��&$ՈP>��]^~>��B��]ud�RPb&3���ʃf�r��믲ͳq�@y�Gߑ#//y�L�x��ΫK�矅��)�x��e��OWPo���Y�<�6kҊ+�T�05s[ĔC��%�8��2(�q���엜���+��7,�.2��"C�c�	��i��aԉ��lĥ��m���@� ���Ʌ�9��"O��y�(���W!~��^8��*#��v�|2�'Ɍ��c�lp����^�]�1VTÒǏ�3-�^�����4l'+��z۞H�*F&�����y��[ ��?�Kۘ/lW@5����/�%��"&�\Z�)�F$�0SK��Fa��;��|��Jk���Jˆ'.����m�y�{�Đ���
����
,)��A g8�7vj�Pd�E��
�Ś|J�4��%_節po*'eަr\���O��^���n���vJ��E�!�������3����/��!=�`�䝣fOǳ�~���M��~!Msm�������Vw����1��I�H�+�ӗ����!�lf#����lGb�R������;[}«*���|gzb�f�D�\�8N/������W�Ul��6�{r?]Ho�^L��-b���h�3�}L�)U�"�y�e�!��y}�^5qs��t-S	�P�R�_ݢETA��N��!J������-�5'��C	���A*w�0�/_.$�~��t��$�{	5��_h��2��*�`b�`+��������{��B�};U?��u��I�?q;���;žnAς�2]21��TY2�>ݯ�r�S7��i�amj��n#�Vrw�]K��CB�V�
��?@f�&�ª`�N�H�C6q͗av��ʋ�y�޹��1Vo%�!��.fMz�A*��C-X���5�s&�򘰃S�Vg���@�W�h~�Z��0���R>!n�7p��Ҝ�������8��u��Vèē$����N�$�G�ZN�Z-y,�
�<���xҤ��V�h�~�Ѕ�
���+��j^���EW6ӝ=��Vq���pΔ��Sl�����Kk~���A��G�����f�k^�R,pn�{��]���~�Dfk�f|�����Q�!t66߿}38n���Հ;սT� <ퟳjZ����͹-�:2]`����I](�Ӌ�;�[]�&JI8�/���Ru钗��w�\�"��Ɲ/rڮr�vl�,��:K��U�v��]��x_u��Y8`�S�P���Y3��k�"�����Q���=\�y���W�^�Z��͛)K-�{ss�1t�t�˘�<D��^�M-e�D�ޠ[��C������*D׊}�:;KR�,�A������y����?F-v����v'�[�����
*A�7�������[�7r'��c�W��nJ�k���ț끝�xz蘺�����E��`]J��r'r3�
�%�K/GŇEU�6&�}!~q��O�����T-�!�J��V�5�=��w��	#����Vw��)܈>�]Nچm���I�P�L(�!��~�k��ǖ�_{V�j���Ʉ1�ġQ��՜��uo����(��_o'��(�o��!������dz-m�1�ܩ������8������-�z��Q�4Zo�(C�[����S�df��r1X*)�2m��E�=3Q0Z��.ç�É��[�����@X�k���^�C���>��ͮ�,�L饫ܧ���.o��ܺ��ݳ�Dݲ��T����KV�!�?+  ��;Ԝ��B񃀬���Y�$GI�T��nDUʱa<}Bo����N�������B@����+��kΕfD��d��&u6�n�Ú���t�i,��a��Y�rKrf���h���;+����*�H`x[�Ҝ;t�v��M���d�U��~��/-#��p�?.�F�b������Ǟ��tD�:� n��ûIo��%��B6<�BǢ�2�������"|����sڋJg+껭�f~���>db��8Ԥ���5?����� -��,����5�~8�����U�*�@�pvE�Z���&���r!T�	
��=��e8��4]�,xp�Y1�v$�3 ����Lu?�Lz̀�V�@����n��C�?i��`���U��_���>�t��%u�����z�3�]
!8�ԣ�n�N�������h+�	��nJ���u�:������Pd�-g�潠��H�3������5Ss*�����n��ƫFY!J��&>q��_�Ή��DHρ���,�L�;�x$~�[D�rQe���*�WZ��DM�٠6�Cb��g%�'��mz�9~�̫w2���=r� ��@<ҪO�5+��X�s�]˹������^}�-��1Q�� ��F�¯߬02�sס��7Z��`�m?��ǥ�ec�0P׀�J�#F��~ W=]=��_Z	ۻ/a���&�9�3�1uI���co >=�OS��[�Q�8R�Rt--J��O�&��51r�M�<�x}	������:�::���Kk�7�n_�N[c�:'g��^�����Nx���#����̯�:sUE��E��fxSP���Tl1�z�o�&�cN�9�ϊ��5���(��@k|�,SV���z0-�E��ڴe��{�ցM�S�L)A��� gY��YW��A��x�oK�mT0^���tm�S
���TF�����j,d�=�,vNO��;���ev��n����=N�٫;�O[>c5<:��4�6I@Dc>������=��i]O�I*��k���^��g�$f�<H��7�ţ���k�p�u��do��Z����C��_�$u��M|��z��ں¶(I@$��������t4����_�2�C�n�6&eifSXxEw���ţQ�s�'<o&��P(��v��EU+r�R���hk�S�\jj�ă�����K�8�9��=���/<�T4N��觹�`�r	��w��g��z����x~�ƘITJ\�Y�u��UΎU:	����;(g��3�yp�oW7S�!t0H�MCV;��:�I3�d�ގQ�	�����@-�[m�=^�K�t��]?���|h����h��^�5� L�G\yj��@�9T%�x���h�"��մ�^�~�N��:A�.�f4����V>����|��� ̶2��fZ5`����7�L鬶1���l���k����▦eH[���Nl���}�S�ϯ0�[S��H��s;�?ޢ{�T�xR����.��i�����L���G�A�sf��S�y�)���<�+�%�K��2��SK�bU��:mr��9Az�Ĩ\�v�D�'�pu��2��O�{"�����*��?���,�_K�}���p�����Z?,����(�k��nX�����7&�4���}&�=�UQV]f��2�::�#w���7���F���b��K��-bI��]0��5���؄��_��E�7~:j��b��T��F����;b tЌc$���B�@NT(0�Ժ�����1�ȣYVO�I-����3�Y�T7��h��b���)�k5�b'�h��-�bxɬ��F�ej�c����:�3�Ò5Ġ.�bu$�ы�>���I¾���X�0�U��-�*|��\����F����1��W���6�;{&:kx�Eh�%�pS's{PfP�Ab�~c�%ᰅ3'��L���
�<��[�ܕ��h�|w��A��3WE$�hъd��J�����G��.�n5���9|���ڐ!�9G�I�ַ��J��VQ$���li�4��*/����Ţ�;;+�F��CR�|��I��>��N�V�^���f�V{f��@Ic�ե����	�b��0�G��/��]�>42V��,T��$u>l,N�Q�wlԬbX�����b��
�Q!�TA�!�)��l�����_v�K�R�K
��Ҡ�'���Q�����0͑ք�+���Yu	�����k)Ѭ�L��7
q�/�%Po�b��pޮ~�]>)��Q��G�e��a�-q��̗��yKg�'{�����y��޳��6���x�-I���{�BKO�3J:r-b^6}9�2~A�DȕZJ��M}�2�z�D�V�@��4�� r���ǒ�3kn�w�\�,R'1O�&������p ���M�Q��_|ݧ��=#h�#�xT����i͙�4|3J!�v��m�ld��}W=��PG�U;p$jΐF���o�c��<�+�<vF<�g?f�U��<}�-ҋ���h�)�t[�����'S{y�1��~���XZ"Y@N�������Ѱ�	T��,]\��ᑉ+��x|wZ'<L�e�\!�/���H��D	6:>�Xy��J3`W�4�yK"L~
N�2ڼ�1�Im�5�!�\��o۵�"�_3�n-���NK��f�y��5:X�v�RfC�;��t?7�=��Z�O;���UP���.(��=k}Q��B�Q�V@
$����M���q����@�� ��+�f`���N��;<�6�r��W�����g��	<�7�hUkIf*4�}����Q/��?�X-UKs�d0��XB[	�h�՚�v�Q�֭�^���r���2p@��y�߮��MR۠��J��*�Xs��ꎅ���T�nB
x�]֣|�>%�.��ˋ�·�g �¢�_��~�k��ܯh�O[�������T��?����J��\��@f���ʹ��Z��2lV�z�s��b�H� �t���p�f�_��!��ٓ5�Y�-�� .�,p�D@��.~�(�ͦ�:�豈C�k��x9�d�J��&}D!ҭ��k1Z���{@|zf+����?�`L���A0�ZR���/�gO���U�&%�M2)�Zc��~�| �mjݕ�%�_'K�P�7f�y 㬐���z&B�^^:)x��O>H��cƼ�}Tgʍr��v�+� ���Ǘ�à�NQ;W��@��'�r�U��a����� ��@��j�_H��A5=qm������0�>�5���P�v�jg��]�Yb�2ا=���l#,�5�e�O��牿w�N;S�/V�GF�����]�t�?H���`��9��j�%,����p��Ǔ8Ju�{�ފ,�
I�*��_��x]I;�e�N�k��Qa���6�-mDX(s��8���"��_:{n���C�b��c�c�#�}p&R6m��n�?q�\Զd��r+e(��������7������e`����?7�D������n���4���X�t�0m��;�«�9�rcL��f"�ٸ-5�[O/a��[�x��Y\�K���v��� zh���`r�I�jE���5+�J��F"���L�n3�3hJ��ՈUFA-L�4+�+=�.�H�a�w�,bWѧ��4r%!��L�e�_օUmQ�x���Z�eJ�yQ�&��� 0�Y¦1-��c���}�DW���"����Q�t�_{���
���w��_�z��������?)�I��N�ԛ�]Q��1)�J͂+A��l$J���2/��Y�:aԷ�?�Z�^�u	��Q�X	���ޣ���0{����,���W��E�������7+J�A�t�ǩ�����=��s�;��ܳ3���>�� ��n�(<�҉I�}�D�E��Wiۿ�@����z���t��Jd;q�\U���;_�`��	L�����$*�]�c�Z�(��T���Rg�F� �3� �	tͺ�2�Pan��$I��f�յ�V.���xF_nuMu��x�J���z[�>\�~���t���ڳ��(@K}ap���t�1��=l�# )�S��D?���GfdD!�p:�!������c�	��F�����
�C���w.�:K�?��Q�_���-���@�n1Շ����|�7��B�*�q����S��D^��g��.�ڗ8e���QP?�?������sw��del��;B�va��˄w鐐�8�z���/E#�'�;�y�V��e����
�����]�pF�a�qq��{�PH�n#��O�f2���������D��˽�rv��6ui�ěն��,;~� ��E{��0Xx���ѷ�� &�K%��Vh�G�ZR�9c����s�qAZT�0� �0v�+��P;�=���D��~5����MP�@��;�<��0�]���'������9ҧ�:r��d�d�yO��F�3n`L	�k���\�YI6���+��9|��;]�^%P�1B���OT`��f��x *q0��TZu.�ڸ ,�R�*���3U0������'��%I�[ߏX�4k�$[��V"�9��桘��j��s=i@��ǁO����QB�m|�"󡼊GD�@�ʶ�09ɿ�,�W�z�+�a
�d����ы^��_�P��'�`5R��͓v)ɛsiR�.�.h-J�r#{	�4>��f��I�	���VQ�^C��V.Qi���ߔ�5T�d�l�TiM�<
��(��6�P���vC$�K�@��$���[w��[d� @�2+%[-�����4-�ܘF�-�	-È�C��&:�JVr8�P%�����ϻmOܽJ'���	�Qx�~]��^?��(
}BT�j���<�'lB��/�����s�;ؿUǬ�b6sa�!-�*֌��2����$�y������<����r�,\z���$����g��81K�ҋ�r׎�Lw2�����֯�_e|�9�L�9��߆����#"L��;	yQ��s.Y�&})��@{v�5(�1\���%H+W�8e�ܠm�DO���p#z��JQk%�9snd���is�JF�+�1
@6��<|��b�zbiUh��n��!�-8d|�0e�fX|v���!��h���0Mo��A=�����:�M0h�HŜ=�sT/ڒ��+~֯�D�N�w��c��H�y�{S��N��n��b2��n��t����Z�ߘ��5��q[�����Q,һ����t9�o����i�$�r.)�b&sGz<�Q���u��E�}7]��Z���n�z��t�=��l
����F6U�n��|M@N���/ci�}'�0V����[����H�/��Ň�,e�(��:q�D(8q�{���֗�
x�8D:���W��z78��u����jɅ^5�*��XP6�0�EYZro���s�!���O�!Q�7�F�}��]=
)35"���[����c��TjӉg90�5^wi��ɍ%�l�=V�(�����n�V9|�kcV˨��@�ӽj�l�NC�u 7h��tc��7 �{��~U�]�N|-L:�b�!�����N#\j+��]5V1��� �58�W���*n"po-TX�k��0���	}�CYSs=���{i��n� �^=�F<{��cu�]��C���y��RXZ���=m����Նx´&�W�%e�$y��,��f
��i��ߴ\P�����x��V��;3�'���Fd1�K��S�����"�֎�r,�4#���>��2n ��d6�^Q�X�4���F�%��;�lD(�dx�
@���ك���̧q�ݔ���Π��:��d�Xӽ���r��7'�^�.��c��bw���[�>��Օ�1���jS�Vyt��d��+q�'�k>���u;�"��|/�;��:�x�y� ���I��[Y�t5��T/�,���h#����j���]�$���Q|�ލ�p��_H~��.qKc������꿔!>���8��k�宑��B��z���p��;I&B���Oƫ)'�`bW\�I*���lqp����B��݄�I�t"!ҮIm�2ElSw}M�µ8^u+��9���c�g��żE��_�p�&�%��>9a�"s~����&�E�N$��Nb�y�H���[g65S��׏f��ay�?,4�;�v��R��8������f�?��y��p�18��CHIڌ�K!)IQ��٨�#A_��x�  ����W�y��-�@/���g)*Ħ�����X�[���|�e�6��<�'���K@����9}U�y֥A������o[v�@b]& �4�7�t6��%�J�VǏጢ-)�I}���I��
E��҈N���ER�36n�˂��1�O�k7�n�C�rl�[�O:sor��N��|��/��\����1��=��ae&���lT��dB�kn�xu�Z�֑�����ևΟ?���Rn+L;�~��|%�g��haR�����YޑcX�ՎZ�ތ�U��G�*%�&��2�t��O��]�R^�.õ�iĮ~�A|Kd�A�ELlgq̣t���aլ>z�8�ϸ�ۅ}b��1(ٍ����n��z��!%Ɵ���44�ª���C��Y�&0�w��O�x���[�q$�����	��L{��>��4�.Hu���hw�jl2?��~����������S LwN������z�3��Zyc�Y55������Ͻ1x~���)��֩���ǯg&�A^��P_O�7�vFR�ۚ�����]mm�>��b� l�G�rHj����\QW(���zBM�l�pJy�5�!B%k+��F�>?�26�r��Y�y����m��]�]忉��Y�}�8�(-I~���cM$�j��v�C����?Я`^��Z�Xa(

.�E7�'��Mg�bO��l��TVGʪ��v ���A�k"B�2*ݐv�0��-h�\�K{{2%���:l��,�_���8�[�������D�9����S���*d7���3s�06a�&���2	vN�2�}�Wj������Ko�"9q��zB;/<w�����+jG�<P#V���i�c)�;fU���~��x<�"�55Ҩ����ֵP�#����DRQe)�`L3��������"z�{���U���O1yT��i����T��oO����zRA���
;$�\Q�.4"
%���]�p�oԹ�&�/�DHW�\G^׽×����'�7h�1�{�H�D�����Y�FJ�Z�1���)�M�l�j�Q�fM�J�v��ײx�~㝎ÓP��T�ED�Z�&1 �W�79'o�:�[���f��+�D��D1���D�"y�_��7lH�nc���b5s�^��6�L��&j�i�3�M6v�}߅���@�ټ%ͼo�PU,?�WR���~e��Al��B��nE_��.�	�`���Ԧ[�ӎ�Ę���<^g&w�
	~|�HG��^[�t�T	�7~^�ȱv$ol��ӝ��K��s��H�߾��ѯ7s����l�{Y�i��	u5�[��$�M�
��X�I��� ����V�J�5`Υ�~}��,�/Ԍ �k4�X�����}5���5����3e��.p^7l����� �=[��R
#��(X�AQ�<��il"��l״�Q�f���53}�	��}-�R,���M�:�.n|p�N-�}�j"V���U�*E��b�!�린��k���
Q��3au�5�L_5��q8[�0�fm��E}�A�kԟ6�����F�wz{K��U�W��'wKa���?|<���v)'�� ��y��H�\`�����G4�$F�8�0�λ��ƞ���D��dק>XP���V�R��!>j�h;P�1r��b@�lYŷ�m!'/i?�
�;t����{9�a�V�Ĺ}��}��bA	roҾ3,��D���d�"-��ͅv]6��ࡢ�3X�eD{	��$�>�A��$[~�6��auT(Ȯ{��R@����X��$P����T�����.���3?�J~�+�����P�۩���;��6a{Kj}�z��h�Y�^w5�bu��[wht�"&#.�q��U��{���=p�Z�[�nw{�L�v�����n3�aS.S�r�����]n�b��+ ͬu(_���U������z�l�	�^��婖U6�H�k�k�4�U3b�A��-?-Y`-Ź�W�Lv�9</z�U\�7�ұh��s~p\����q�C㻌��xڢ�:�-�����$�9n�)?����w���P&b��Xܜ��W��~�W�p��RCcI=Uс��,.k�/�`�&/}��+V�(:���/�0��(���2Q��˜Ẉ�W.�sY�Y��o��1�{����pw�`���,���9���w)!G#��S�诖Ț�C�M��b&��lntO�(�-0�#�y�2�6��=p�X_q��Q�2��y�p��[�����p6��e�_��P)I�C����(��iyV����v�b66g�;�Uu'����܋A����9���=��S���_>�m�>g����p�'��������#�u�H�P[�47ͭA�}y\��P�7�,M��l���^���h�O-�2�Pq���ءR�V_�~�l�촒�
�����^H�߬�Qf�l���t��7��x�������-'{sjO����p��
7+N�2�h�N���=�!k9��d��_L ze}��>y�v���3�^�.(׷��2
�_LE�7B� ����M��D���9��[�>����0g����p�L�%YNF~5�|G��}�����L�&y�S����Lq�n�Q
�;�_������3�c�����Ra�g*����痢��Z=|�a���ߘj�Cx��F$e�g�=�J����R��`M_��j.=2��}^u���Z�l�\h����/`R4QV�|^]�V����7�f߱���)���X���E��P\�U�������i?�������mzO���%\��g�}?
�t��*nI��~��mw��f�����}Ew-��s{��_���̉�GS+�*�l9�"�T�u�R.b��3ኸW`*��b��9�����Ь��;/z���|�,ɌH�z ��h�NӠh��*P}�zs���D���0ꊸ�Q�990A�=�'`��ͤ����f��;����-��^iݳ��"��mţ��A�r�Xa4�8��TX:�AH9uHxX�m� .�z�0�
� !�)���{���h�FNW;2���C�fWv��g��+�L���z�|�ι��ZWl�j��C0��	�m���m, �<�n�8+��G����0�>��QI�#�L���w�oᠫI((��m�6�ʧ �iziU���]Q�����w#%�&�i.kӓb��ݳ��\;�$>}=���y��b2����v�t�ܫ)s���j��u/B���71^�y w3Y��ңu����x���e/����0P�aL2��݈4'�"�&��_i�VRy���FB�Y�)����{3%�hH�k}��Bc3�K{Uk���K��5�D�t2̴"Q�BG�h���Z�g-A��.���IڛU-K����'S�=��i�SK���?]K*�'�9���\Q�/��/��걠��;<㮎WdU>�8Y
�a�>X;&K��y^"I����%ϓE�#��7�-��͡����[W�ٗ�Lr.���|ľ0��~g���䊫���Q�e�T��}'�+N0��θ.�V����3QV���Ʈ��TZmE�jWì�㠾3I�0���US���S`�c�#�r��J!�b�sQ�������kJ����������՜g����CՒG�W�h12���g.�صv{�sN� ��y�8�#����r�J�pM *�[C����{pk���j���*���F8�d��l�!��>�ij	�]�����US�,%����$8�1.��&��%ndD�U3��f�]�?L�eX[��=L��ZܡPŊk�b���)��@��@qwww/��,�����y?���~�̞=���:g�pfis��ik���ؼ��9l�f�M�5���>�DJl.���Pu��0s���{^[�P��O>�������[�R���c�*�����O�wͻŠ4�����*@��c�PV�^p�h)p��7 w*op�{r28�&�D�
 ~%�QЙvĽ���I0�4�OZԸҀ�����~��W�j��x�X�^s�ho����v3@�B;D&)տ�������K//���_�;։v�%��z��K��j����9����vz���"�%i�O��%_=1C	�<��:J���	Kqׁ�z��V�D�����2v��}���G�:�y���O�՟t:~7h�U4)�%-�+��Q����*o����=*݊v�e������a���'����ؑX����{�%�Q��������yB@xm���PN�W0�r�#_X��V.��26�1�iF�*S�aR��P�p�}�6=������0h�-�]��Y� �.�0�Q$��հ��z0��`�x�A`����uP�����5Of�"줽a��0�{��'�7?����G\��ʯ#�\F�v[�1��S���	�r�裾KҾ��(jJ�m���y�� ��\���V����G׎�*h3�\�c�$��ċU�B�¡�V?��f����?�ٛ`ɮ�v����=����0Q��3���g.�|���>���owVԼY�	,�ɝ�������bZ6��Ɍ�l���ć��}pL���X=�R�Vim��ƿ�7y�๗s����w�Sv�V���W�I�Ү��d�F�Z=�Jem�􊷯.4�ߓwWi��al{�Q8d�YS�?:��"ze!	����iQ���X���;��_W��X�9h<8Ϋ���R���Q�����L ��p/�Yg�a
�LB?��E=6��U�Ir�j�<�n�>xv�*�=}��qq��<D��ϕ��R'z��7����Wm+R�};��)}.U�x��	�}M��yr�,��ȉ��VF�-@+��~G@`���o�6�R)�T��vL��.>.�����=b���]Q�7�ͭPgI?�֔`�wv�~�������͘����O吸�cgd*���X�Am��q^6�ҳ�S ��s/i�	Be�)�����x�~�KY�c�ňi{����m�����i�[�f��b=S�}���W�/O�2+@�F�6���Np������q�BH2��Cx?�|XY�{T����;����h�zF�fњ�QZ�Պ��H0%PΠ۹5�{,!�z�2�cβ��l�CXɿLA�&�y�I} ��.gS�-��x9�$�d�*ipp���v9��{R�T<1�Ll����:0���HW|� ��ʦw��Y1z 	�{Rֲ��}|���Ӝ��m�|�,�ٵ�(�T�-����ACMY����'m��g%,F�N?��Q��@4a����K�D]w��a����3���l�	��:�ևhB=���g��3��6e
v�����fO�p����=��S��_�^�/Tn|�Q!�va�8ˮ�M"��>/xj�]�P���n�a��<�рO��`���&21��Պ2	����͂1��u��@G?�V���sR�
��+ʎc��ϥ����V�?h-�v �l�o��J^ףB:z}lhU� 22�u�W�?ā���������=�I��}�����-R�ysWL���xd˼�:�_��&_;y�|A�#_��^���p
̯w���DH�=Ie���#�(˰U���%�a��X�+Y5,	�]Z������p�O�����n �«ء��3�o��w�n��rڋj�4�8hN�7��m(;�� �#��ds�wm1��)�'1A��E�*���d7gc7F��x}
����ҽ�K����.�� �������	��(�HT ���?6�Ծ��0B��:���S���6����oz�3Zs�M<�t��q'�:��DV�!� �HQ��*xw��撺���v�)���zU���2ԑّTS���
&�L��Z����[��U��`��n 嬣��"���o��nǀՉ�yT���6Vm�T��`\�93��o)y�m�jx�L~D������H�rv��tlv"���j�Ι�BL=�i������0P�9��`c>�9:\,Ϋ����}���r����h3���Ȫ���w=U ��?͉���P��R,U"�b��&�$���77�9�l��m�f�b����M��B�Ϋ�Gzz����#:د�[R����Hi����n����D���=W���b�e���8�vR�qw=Ľ�fz�iӶ�!���m�%�B�Q�:����@8��uC�g-����xfWj+�2��W��Ÿ
Nj���:��\�O6���]7�����U�]���*��o2^5帙C&(JE��%�	JF�g�vb6�Wy�������&~���#y%�..K��/�c����f��WdQ���A=Ʉk��~��يn�_��D�t(�W�
�{R�Z��
��:q���3�H(E�I�>�VV�X���:Wm�1���}��0���/}�ǟ��e�?8��X��'�xpaBN�w>���6,�l��z'_���� �QC�Q�k�y���޸j�_DV/}B�7+�@�/n	r|�B�1
+���s�-��- ��O��Ujo��Giu:�t�Z�����S�T�gn���n�`�^o�ڨ��u��7Hc�p) �F9��)�S��wr(Ոn<�����K���bGD��GK�G�2��O|y'򿷏C�.���#��WZR����^S$��b�F����:�̬�A&�@g�3�[+П
�/i� �T���t�.�O��<<²3s��7���C��cd�},�)e�n4�Мhc������;8կ����(���a��فq����;�tIZb$0�����d3+�-4@�Q�sD���[s��,��Rr�]�p��5��7?����](�$�zlq���J#sB*q��%CY�!�7���S}��P��!�b�*I��96��nM��D����Յ�gO@d�.����?��d�\�ϽT^E�͇_e�I�&��-�x�%�/����O�S��Ku��:ҁ#k��mxM��g�5W�i���C�{���go]�mN_���~\Ŧ�ҙ˝[��������2E嬑b����w���5���*���[�f��"ޣ��>>���x�M��Rh�4�I0,�m�\�L�|����h��Z���u���#���b�ʜ�|L�zE��H�>'���r�y��Vv�a�8�_�k8��L'��b �g�4��v��3���9t{H6��)�K,�H��J��u�!HjT�`��1W�����N��<
h����n��ө8��t���4W�e�J��B�	45�z_�૷�<�8a&؋Al����7H�AM�v�CH����;�[���N.���IE'�S��3-Y�I�/0\=@�ˇ��2v�w��gH��f���O��Y� Z~\�2 U�fid�31;��^W;����@_��4�~��#Sm���|��ED�����˿���˯�6�Q�D�A~2�\��Nk����`a����mv��F:U�ˍ��U9~�� [�D����hj�p,А2U�V0)�^BL'�#ar�ܡz��H���N�|f��^cC`�0w�Z��:ݝQ����=A1<9~�}��)l�9l�f�2a���Dْ��pڨ� �Ȁ��A��(Z����\*�i!�J+��l@�^>y0vl�pT��/�,�B|w-jCO�v�yެ��V��؋u+�Ϲ��ސ��l<?�jU46=n���sm�\�lO؎5n��]�[�Ӛ oʌ�����v*��3�glG%���!��X���tc��S��,$����u*y-kUawg3-�����q����:�A���r0�Vt9ֹ&��XK[u�{�����na���V���BȔ �10z��r���Os�t%���軇 T=�A�!Pr�ߡ�C<�V�鴂��^�8>u\V�2�@d'�9��P����p/#r��������tL?-�0b�����m�嚽�;����^��D@Afϋ�w���q�;��|��n�5=�?�z��X$["�/Z�����p���G��J`�Vr����S�����;�2'�=�/��˺�׭����i
)��-2y���{��
����
��o��L�>
�pf�Y:ô�n8!�g<�B�-�
[�G��5�Ȟ[-)�[ma��}���u_�j�;�x�$�2�U�tK�N'Ȯ�'q�tQ%K�e�=A�����0y�a�;���j�����Oߔx�`&e^��D����f�>��qhp��&��k�`��"E��98|J'����E� ���Ѿ%G[�HS�*?a�i/�17� �Q�#��J�m��.�W�)�H�pᾮ; ��+|Uk��ūU&���9YdYx뒀C����z� �B��-�Ō5�iv!7Z�俣I���k.�<�).7UVk�q~'{���"�<d��ג˵obԿ���<=$#Y8���Z�Tο���R�����:�Λy�q��hy��3���o�o�����C�<BB����S}��ҭ"���ǖ	�07�r!�#ƈ]`�U��,�X�VlB�cö
fx���!j��ԯ�E��~i����/�ft�\_��$� �U,���5y�I
��vn  �o������u�w�g�J=)Y�Km���OH�t�7!H/	����;l�x��<��k��%^�?\���(N�����~����>!ONN���6mx���}Gm��x���lB�	�"k��,y�VW���A���7��W���.yݕYyzz��񹝞��5� b������=g�G����*9஍_9��2_�px	�VY[[]Cc@��|X�1�AT$=�Z9�ù��{�ɛ��W�����)���ϐ�J�;���\�ᔛ�_t������ߐP�kċ��맃�ߏ�:=!_��x�F�\LƑ��b�©���8 ��%���i<�L�
����)����6.���4��۳!�C��Ft������Ķ�sqK��	�k~��Ƃvy��o�ci1�cf��a�=����������Apz���qc>�S������E<��Śu�Y�^6�t.��v��l#_��7����@5�'�벓����{r�-�ˢ눔l��������T��� B�rBE�5��hl�/TNY�ߒ����@�ϟ�R��oHHd�ٰH>�f8��qK쳓��fLVc���oV�����&
��鋺��W4�̞]ѧ��d�����(�9﷈���f�?I�=v�6��"���Vn^;6��4�k���U���AU����_���.$����\Y�oCE���>��f��!������'�]�7��K��kj_^�]�c��3l�U�5�J�ք�6r-����+���ʒۆk�N�q��ʆ�����Ց�kY�su�����@tL����a�U(�D�M�ET�\(0�� ����r�w��AXH(<[Ľ�������<����q������Ъ:�'�U��/ZNt 9�9��:���[m���K��1�����@a���E9�\c�ke��'B�3A��
��A^��mw�MzTs����؛ᒾ-�ϱ!�L`��üR�n�(�����J���%1�����2Ah��9�[�������$l�t�4��8ZJ��5q��Z�B䢺�(4��&�j���gH�����x�<��elEo�Ae;��&-J{�����/�\XZ�'�9���T���=������p��EppӾyt0��7��xR�ןOw]J��p��i#`���َ��d��c%�议D�a��v�Xe������ֵT;�1�k�&����CM������"k��b�t�lK����CF��ϝ�M6ǌ�SKKeˇ��Z�A;J1y�3��	��|���B"RR��F��g�7��*J��]J#�!"*�$$�W��b�iN���vy&�V\�iE |��ݯp��35�Â����Er��Ƙ:AD��`�����#3�b�s\�ݳOR��_-���sJ���w�.��	xAX%��4fg>���L�ؿ���qbhg�� �ڳ��V����;��ӷѷp�W<�eju���ߥ���|:,���tr�~���E��_@���Yɧ#��P���8=�Ĉ���%[G�3�>������(��9�$�F *�r����Z����e�k<����yL�a��2���6}�h�X%�2z���X��>�##�o�H�#i�9�?h�)�џرɂP|���0sj~�ե�����[8�}��.�,k&MC�I�z�8�ļy�l��?\����a�S�����2��)zh����L�x�!Yܚr�5e*|L)U�����]�1c�p���SgX��4!��� ���@N�(�t�N�2���B���O y&�!`m4.L������K��W��4�F����Oi~؊��76�Z/��2 Q�c��sp���M���w��9�o�)���1���ؼ���aE�#Sf��J����-�9`9jv� wr� �-��kj�Qt���H��f,uy4�m#��\�L�P�l�S�S:�&�➏�Z?��n���� ���~Cw����~UI� ^^^�e�����!��Z����W!�_��*�؇���:I*���.�V��Q�*�n\`�(��x�SLS-���^3��V�%�f�L�(=�Z���w��L��[�����C��.YI9Q�ׄ�`%+�OH��K6���X�G���Ә�'��u����F���'W��t7����t�����Or,�F�Lo�������T���d٤4�ǘ�6'G+��l�  ���2~B7"@.�Z���sߑ�3�Yv'��L���5����:r㴒��`��u_G7��x/V �0F��ǋ�7^�G>X�7h�p�jl�@k��Mͣ�,T����@u	�ϳa�Wy\��B��J�����-���
:|�	Y����k;��ڠ�ց� ���Dt���r�Z����<��3�� Q��bL]r��0��9�6�q�Y}���O=��gr3��w?�����qE�p|]ok����@Փ�+�	�,4o&(��>֥k*]`݅�d�����XH*��3�52DX^�1��v|I{,9�F�� ��g��G��S�	�m5����8XѬ�Tws�.��w�?��οa� o��:����3c՞�j��6���G��3�zb�g��_a`A�џw�ǙR�f��2��w+�S�C�*6"���x�rn!g]It��|�`��Z%ژꌓ��Ť�L�,:I�����|��70�j�y�g�p(��ɠ��<����u%��c{�3,��ǹ���	o`t2��>nq�e�kg��҆�_�i��.3e����ՅWa{�]�*^�����Gѩ�������Qo��P���t~��Y�qZ{R[��C��ߖ�x���Y��]���م𗴁ԅ��r���6�8�3����595cB�|?|��5�?'Z�|h�1��Ύ�ujyU�'�x�A�o��u�"�آ�P$�`�#�g�Pً���?���s�. �C ��,���Z�SnG��-wWI�����KQ]/J������?�#2Xn}2е�*���v�L(5��N��	ZLKm缿�;C�-'|l'x ve�l2�͹����H���k��ʏw�Esd�8�
�Lb���nC�ޮ�V:DO�E��cΤ�N�P��z��gXz oy��wBP�<��79&h3\^TT`��.����4^ϯ��#�G�x�
��d��S䥳�K�o� � ��.|v� �*^FM��G�>^��60�@��J�[j�f�P�t�����r�:��f{bB=� ;��_�2`������iC��?��.n�(��!�m�e�;�2�6���~N�I�-�F�I��s��M�TT|W�Z3��;2�	+R�H���>J�h_-�-$��!��#,� ��YL�i��SM��a�K�o�Lo�W^�,��;�{\E���(X�]���\�h.�&>��u�ߊX��� ���P:�m,��X�c�D���6/�Y�Q�P�g�(W6rd��`zלA��&ϧ�۷z���Ռ���������rlK2=� �W$�m(B�eŚ�u]�$�{�ɷ�1H���&`P�ju(
�^O$1�2r������'&�wk�Q�Űa�p<G����{���!��D�ݝ������Ʀ�z�*���GNQ��H��7�+jf��ݬ�g(bơ����c���2�I�j�+X�"M��T��iZ\6:1�B)�&]ӻae�7�rp{��)`����ԯ�t��`o��A+s��ށU�?��R?لa��vh�d` �R���˘�O#��-@X�Z�d�/��� E��s�[B����F޶7�W�ӗ�/�Ae?�nb�w�eZm}�ک����[������^�}P��s��N	Su�4��za�p=�UMl�Y_Ϟ��J6��n0�������	[�����h����J�w�ǥ��z&A.�B�gp�n�����*?�mU~�^M�q̲���#��/�0�$�]��`~���-�S���u#�z��P�T���P�*vyp$��GhQв%r%}�|�S�Yj�j=%^I#a�!�8��A.�eE� H[J���E�'�{#�h�B�t�J�<������6���8��HB��˫+u��=���+��.q��F"���P؁b�W3��X�Ek����}�W�Y���Y�_���N:|"��񅨟򆛑�iY�@��˫�DU�ޞM�+��X��d��y���"}�{��Q��Մ��3�A>�!����)�˻������O?�:�ޛ�m4^����;��f�O�;o�^d�����UY�/&�7�]�K];���b��Vy�B3��)�0sPD��@!b4Ss���N RS�+���Ԯf���!��g�&cQZ��]��<��ʴq��g������?{x/6"��8&����Ok��ӾUYE��\2����J9��2�"s���d⭇�L:���`"6�4O�ۘ� �K!j��;F��j�p�΅�\�d�ܹ5q��9�=�Q�*+�q���,��+��&YQV]�nd��x�5v��[�R��W���d�L	Ua��&��3
�M�.�6�4�ܫ�,[�&�
��@k�I�a�OƧ'��>���[CI��Me����[V���~�������r+]Ey:��|:���l�@u���4����'���Hp�p�`7��:J��u�_N?#����y0D�>�����Ų�,F����i16�%��6�� �Tr5��<
q�^�����wp������R�Vf�q�"�oτ�/�z��Hp��̴wI����.��_���ӵF������"1�v��Z#��Le
�$��!���ݤ����f�Q���ѳ����	f*�u���Ht(Vm�~�˗�b-�Q�*��Hh<5��E���6- ��㠕a�S���4�pf�4�e����Ih�Y��3�����I���o��CÜ���F:�O-V�=���$���.��u2zu���;	�����7}V{@����Z`ΙH��dQ�=���*�`�|,�e,cw���CL����
�*��:�t�\�Ȕ��w:�w�E�%�3�R8rW�֖��Z�⋯#ߪht�p��y<r��6A4�l�A�(.�k���n湄x��L��[�psd8�M]����Ȋ�̶$��¨��唡�>�y��/+���ȓ����<]�.,4'�7~�=\�����T�'2܅T>��[���9�Th$�}�o3[2^�� �h�_!�X����8c�$����(`��v�P�,B����+"4�׈Idis��r�;Tg���t�y���I[��z�m)Wu��Z�M��ۥ����(f/�}Ef/)������< �䓠�!_�
4�Jw���&���1�}M����4��䳺��ģ�_M��ޔ-E{�\��#�ʩ�fx��DT:{��!M㾰��ڿ��&u�pg˻�,�G[��^Yw3"�_ON��;i���a(fe����<1ٿΚ~r�:�m����A��{d��y0�Zb�5���=x���X������o�,d���w�Zi\������7���0�x�B�UʖPzO�Fj7x���?�w`��(��/���%f"�K	9�[2��{�h���!�rd�h���&!�т�(��-]ʊ��^`Dh��˹D��U�U�t/����A�X�R��d�w�G���m����&��K���X~���m^�P�
/eA��K����k�x�F�W�.����g��0B�H2y����q����_��ZM�o�Ϻ��ҳ��})?����c�3;ՑN�UDz{w���5�.M��fhx��zwF�V��3�p������KU��%8��Ƶub������_r����~ṟL ��\~�~�c�#�1Ia�~��B�]i��,�[��n�j��am�$ov���Ul_t�oy�s�nZb�Y0b�p1���k��q�,����j��t��[Q�^;�ư]�4�V�'6 &#���� d���I&���@&����h:���}YYYx�Z}['�k�O$6O!�\���RZ���Y�� �>�{�rJ>u5��3���(6����X'e�Af%��J̫��c����6���!T�s�X2`sfy���P�\�?�S*�_��;9��cbk��Լ�A��:�ݦ{KB�j%���W��O���U'_�A�[i]`��{?R���.tc�\Ł��w�:�����l�f�#��5ק���Y�?
�^yd!�J��> �Y�>-8��J��L�1���[�:�yg�m�(L�#~��Ɖ�v
�L������\Z�/sB��������?�3_�+��F"��nRT���{������G��=pDM�()YE�.`A�	�B.��>�&.�1B7w��9��[?xdT��BksF\Re$�����xh�k��I~��� ��v ���=Ykn;����'t��<ji�\���4��s����m� ��p��4QLU>!@�� ���������834?)������QT�l��"i��{����/�q��T��nVy��Ki9�=i�ˤJU��U�gjɷB|�wM�>����ZE����94XA�����5W�~yZ˹��rO^��hX:0w!�"fszQ�-s�Su�p;����Z��w�~�f�,�Ab�-��������Eϭ���]�X%Ա?a.H�@�p�e�ګo�w����Z������/ЇS5��E��oF=AM�q���*Ӭ��Y��w���p�|!�3W���	�r�~b����Z�Oc�#�p�AbV�JM��B)�+Lة-lS�ڔT�A*�s��|��Ej��8 �=����S��^X�-���x��f���<c<��rQS�" ���һ_�Ki�;��8�k�NR2�(��5FZ!����rJYa;���fMv|��^�#'_����0�(Q��pG>�'�kU���fկI����hl�y��X�g�^L��Kt&Tb[PC�[p)�^�֘�-��D˿j�_L��/=8V.�PToW&R����%e|9�m�Z�˗8���u��R�	,JU}�f�e���ψ����^XRԖ��,�H8�guw@�ݠ����5�����p,�|�bb�11)�7��0����NAc�����v���I��T��f��lۣ�g*-�QbOHE�)k�ɯm���W*��/b
��E�3͗�TB�>��\�;�;�^V�E�'D��>��"U�����B��Gr�Ɉ,�Â4=fǍ�/Z���s^���(;�v�H}1���b:�d4�f �JP�}�H7��'�|��@��Bn,�u�����E��s��{��6�0�l�G ~�V��U����d�
���h�#Sm�l�ӿP�f�M���N��ޜF$0�uW����x\Y���n �j���=KU������%����	oTT�T�'�8*{�4��1�>a�"`����O��JP�w� N�lx� ���2/�#E�A1��C�,T�T>�0$2\Dh��!0>ig
��(��\�4߹Ք�7�^������������>5I��
]��0>�并lF���r��Znl��uR��?mL/�FD1̢�R�F%��{si?�P��I}b��)���P��ҽB!��/��������8�DU���z�Z�w#::�(r!�(r�`_����D�F��.�[��:7es&JC}?w��Y���׾^�b�g2����$Djz)2;[]��f��:�kI�x#�]�5�����'��_��] �d���ld@�����F�r�-Bt����|�`������҈��޵������
u⌒3�wf#��%��v�s������U�S�%Z~֯(�7q�a0����V��(�����e4]�u��}����w
1d�\�M"N�#�v�V���2�z{�Z�o^]�:r��#���9b�i�<���i��,��5 �š�Q�ל>l��kaS�~���)*$X���v7<�|���;W������%���D�aԯĎhR?��\{4��.�����%��f!��E�7>	�����޽��FE�Q\�����2���u��W�67� ���N��~\s�����=�{��?�Fpٻ�_!�cEb��r�}�"z�SҢ�g{���|~qq��Z�l����|�w�����(�.f�^���T6
@M�Iܱ�l�H:�,�v��q�N 1}�}\L}N��f���DW�v�Ȭ�&���lg{�ç3�a��D�3�E��p�w=�l5���h�����)<�s^�7B����f��ųA��,oT���t	����E
 �\�78&K�t5n�9褓�m�\UM����D?7��l��I=�o��������~���i�$��")|ׅm����Z��	�X���c�1���$>Ҋ5�Z���z6RK�HKKKs�B��W�Φ��d��߯N��]#���Ԅ5�����P�����w� 顡#�W~Z����^�scC�Hݞ7��\d�O���z�4K�F��+�GsM��j�.�k���)�ǬA�n��К�w���zk��'~z�`YѡFY5\��a���cU�D����������x%/��Z?]E ����2�Ʋ%z�`߿��0����|�����-��oY#�DmϞ�� �֬r�n쪦����M��O�c<�I� o8���C��� ؛��_V�
DK�)��{���؂�S�S>���Ţ&�;�c�ɹ�],�D�ȍ)�o�iA��;���)ce�(���[hrN��F'�B�?�V�ٟ4Q�E�Ӻ�ߥ����^7��-D��w���GP��v��\;[�A�'�E ?z�8���c��Jˉ���I� 7 ��.����K��v݊R�a�(jD�a�n��~���{o8��� Y�=���#f)�#c���l�$8h��
��Lڀ����I53_ �8�8�Xv��V�S�~Ee�Զr:n7��n"� �,�J���Ͻ��E��y<h�yPޔ��Zpj���`�����?6[~~���P�`c6�x��t��~����)ֳ���Fx������jU����5􁇵���+�;S�D��,�����*7��`������\k�H+���	����zz�7��`k�"1���gP���ی�o>�F|iB]r�����&�hO�26�X��e%%�kΉOmi|0�?V���+�-�ZGP~�g����;���Q�8���[�9�n&����Q�=����msb���T���"^�\Q�(n=�{瘡�9c� K��Eq�ng�@x�%���*[��7|�t�߫�G��$�..�Z�}�xrl�S���8���#�J�`��6��n��Q�-�h�b����}��"뚅����������2�{����o��J�4��Âg��j�V�$�i�3m�Z˜u�-BX$��s����SO�>zu�B�i�B��*���,f�Y
�������}&Sn�!o�������	�Z#�o��⋗&Ѓs�cX�>�"���2���$%[,�7AWۡt&�O�WPsB���]�=�S���f^E�� q�-�P�Bރ���gUd�����{�Kt.����/q�?Ni��H�]R��Ӓ}@�E�"��9y��� _��-6!����ʶ�c䐨�[Q� ӟOƪ���f�I������.B�]4�ۄZCeQ���A�y��D�8�������f�B�}������r򈑠��<G�9F1K��9���cmF1�E.F�������d�J]��0���8|�-h�h@���(�)3X��%��31G�/�les�t6�R��؃G��eđ�~��S0M�	�~Fd�n��j	Rl����^�.�m�?�ORfA���#~i��"qYc�x���b��5�����9�xu/)M��T̒�=�<3oߵ���
�sm�
o�B&(a�ird�Z�]\�Jf��m .V�%�s��0>Q��+�Z�������")�1q��M�fā݀-��Z���"��E;�R�oi��b�XTw��u@R��|�ǗԹ[yh��%N��rj� .�E�6Pl8�����1(VO҂�Ȋ����Ό4���%#c��%��S[-������������4�e�=Kdd]��[�yZBI׻_���sjp��6��4 �(9�t�� �?�m�R�	�M�7Ab?�,�+��Vs�a�?��?b4v���ٷ_���iV&�Ըߤs�kz��$]�8q���-z����^���c�� ��׈�},��k?�́�	�zo��	�Bu����r� �?�O �.��'#
��-�^�!�h=qb��$tԴ�>	�6�f|r�O4{wF����[@@]},�Ɵ��Q�>��_�TvȗK�1|1�br����i��`��4��v�&�R�!���� �w5E=��s�w4z-���{�j5�O��1���:U��ͅ�s֫��=BV%m��2XM��A��E>o����/����я�F�(�H�D���ՈzO���n/��v�'tf���U�߸���5�zdZa�{��</tV�p�۶_D��r�-VlD���i�v͞V��o�������"�ܔH�Z~t�:}�2�ui:.��o���R�����e�ь5𧻓�8���V��C�q�W�x���7�(q����g
P₍n�`��a�jF�m��7�����M����U%mm�ym����U��ee�5-�Gb@S��2� �	^��Z��b�q��L��a�3��zf��6��37�_!�M�U��@dc�$��f=ʊ]Ji����Br��"X�;�7<���c�T���ثg\�q�gqc߶O����D_�}��Q�x|�z�	D�����~�f���<�5�b�1����~c�Y}��ӽY�X�qA28��m��Yc�=�6��W^*U���Y�Ty%��@\�B&m�_}��4��0�)o�ŀXL�FG�������⻁o���Z<Q�G�'w��k�Z7$u'��V���ޜ��{d��{�T�ZI��-VC�D�4�0��e3FW[P���_���S!��J4`H�Ѯ�A1(�G��Bc��}N�P!�0v(� �2�~�!�;�d¸JS)����E���J�FιG�&�fmt��"��01���7~�
��'���[�OJ��#����э]h]÷����n�����@�ۊD��&����B���h�^6�(5�VC�w@�ju_�rv�u�'��a���M�jS	K�[+?{ d�v��Q?���Mf��:&׫����F{צ�B�&���+�S� F��,o�T9�m2$~�j�pQi���u�Ѐ�J%*J�nCz}&۩�qx��ҭ��r�~��3�гT�)g<<��^�
��������4>�ζjNmsx4��ۧ.V"��3X-���?/���lc�c� {��n���������0��X�&v+�ۼ�����$4�>�Q��\U��� ���a+C)���Bִp4��Ƶ�J61F7��8���E^�fZ?h��J�:�bq�#�
��R�)	���Q�n���YZr2I-�J�1,�������s�0�wuS�B�����
V��:�W�nՖ>��q���W^L��u=m`m��z^?t��8C2^[KZz��K �&0^���t��IF9�M���;�\�z�d&@�Fp�?_6a�	�-�nGO�x����F췳���Y^�:�S���|ݵ'���]Ჵs6�3;���|D)b<fÂS���P\^���iP��U}隝yA���iUy
�/��S$����ԊP�B�4wHg� ��E��z�<�
��nX����(U�Xe�o���A��Hȝ�[��ݥ��UFb ���B�i�঍n�$~���ma�ٮ.e9�WM}s
z9�SSpQ��%���ЏWcC]f⽼s��^~�I�xZ��#�k�,�7�n2͈z������jCi�ƥX�-�B-��)Ŋ��;w�+ŵ-ŝBp-n�%Hp�@p����|�WN������<���!w�FZ�������+>)Ϸ������)��i/��g)L�Ng �1/�,M�Lw LD� ��񝾥r���&�'���rC|Flc���	>fx��
�Wo��.Kہ�6R㟝�D�N�����mH1��x���4�H�vz(�R�*:�TC�����q)70��R�$>�J�а�>��vnS��������<�{ ���pZ�{�a�o�����_�O�%BΥ[��%����a�M�yN@@��3%-�����H���,c]����Sw��p��`�������������N��𕋏��Q��Iuפ]�f����D0b��J�5�:�����Zz��h������*����Q퀃���3mǺ-]B2���v�Z;'�:ϥ��;������%/���5��2��@���q�Zk6Yq��3)�ϬwO�����Il��ґĐ�� O�He�jM5�?[�Z�S�x��=�h8˧���6�m9�%6v�(@!�d[�<�6�faH�c�2F�Ա���d�Ė<mh���MHS�ߏi8Nto�
-��N�_s�0�����!r����U|���'E
�<_���LZ<Na��om�^_� ��YT��$ԟ'��������4A�BP����+_d����t�����f=o�>$�@�`JQ֙7�����-9�xل�:Ԁ��Z �߽�b��L��c�x+��p��p���}e<T �JC��X���-\X����$ds�����F}��z���_�	����9P͎x���O��![�D❽��UT-�3ͅ~�W��ާ��޾�8� w��݅`�y6�jm7��v\	��Tȧ���<�l�A�i"%�(�arƮ�iK�����i��C�S��㿥�	�t/+��[5?p�,�tJ�ϥx>P|t��<�[��=q��`�~���|����<ć4OOg��������K7�'"-^��huu�l�6�8~v���d��!q+C�q~���2��ќ�X�ʥ�u��֟�,�v��m�&r�?V��П�{t^<�s�;, D6ғ,��u��W�}ǣo��wV�y3G6�~�D�`����wHFt��2f��:�En'��fz��I��a:pXFE�wl��\8Ѯ�ƌ�G��Eֺԗ�Y&K!��"2�O�@P�8-��Ӿ��5�?�<B�p�oC@��g�/��9�]S���!��Qgg���՟$�S-f>���(EB���jʮ��p��d|��^{�1�2b�I��)P�	tׁ�H���]�Q�{/X�������N�͛Y����[x�&d~���o8j�{Q�o�DMyx|��݂�b����%<̦�����ޟ�e�A������l=$~�<U��}�O`Ã��n�-���Ԫ]�����VF@c-+�+ŭ��d6�T�y�V���2Mh�UW�{į���6K��J��ᕬJ��Y7h25\���L��s7���]�T� 9L�t0��S����0�=�p,\�����a�E�񽠃��"�Y��D���aB%ja|Ko欲TZ
�R��3;_e�-`����|�o�|�]��,Nm�cK	����Y]� �"G����Y��ԟڑ�z�v�y�<kqu� ��p\ߗ��k� �/�K��D.1�#��n��L-��+gU���8+���v<]���현�� F��K�Ly4uN��e׫a�$��F��i�N*�l�ϣT�7�|�(e�;j��Ռ��3f�C��&BF����D���~���&����ٮ-Z�h��~X��m�]Sc��dkF
ʝ���1_�g��KE���v�7�nnT=u&���.��!��L�Y�W�3�b��chP�$~��80�3j��kOt�dUى;|����}��AHXz��5m-Yq��k�P���߾t	�oq����I|��&�,f��~�zk,G	���7��g���i�v*_�
0�h���ȟӢ'19�Q�����SĠ����/���0y���^PY�M�}2��wVu��*$L���.��~:[9����&{?>Y��������V.��o�ý��o
����9#�#'UC����Ѿ�O�Z�Ѽ�'익�&��=z�d��WMW<�[����hs��L���	OgΙ���{��_�FF��.޽�]��]ց]�h�����Q}�S�71q�|�V����$�
�%�&_�����������<��,:�����7OPZ�nh��ܹ�+�hk63��6�4?���	ui���{���H�u��,�a����@�/0�5�-n���O�����D���=���������'_�2E�vuwݡ4��q|�s/]��l����z�EY9�^h���81xl�\E_U���~�7h��M�ZS���ᾛ�����_3\>{BX��0����V���׬��u���֓�;RD�_� �SG���=�W����)��K�ɜ��g��Z�/䙠�l����/�(�+�����oZ8:չ��v,�%)��fW������ϗ��I��a�U�`�ܒ���`��oQR,�WC�o����[T���6O`��h���0����7�z��l��z�$`�f��9�-�x���0L����fcp�##�R.������:w[}�:���b��1ٳk78%��XI}{����-8���A!��x+v ��~g]	K35�T�|�I��wDS����lIe��f��Mcak|���s���9��h,x�ิ4��8��M{i1D|�Ž���?�Y����M�Y��8S�.��ߢ�dYw}���~|ىǕ�0c[,S.pur��p��n��P��L�>���2g�2Z����������}doE˺wo�NޫU
:9�ۍm��L{f� #��\�0�R�34�����0�r��b�x��S㊃�Al4���i��U���0Dۺm�i��Y���`~�@����$���SgH�&�����o뎘��P]|�*�+�)�\X}i�2^�����/B̶����+F��%�ޘ��D����*5�1��X_�rҬ��V��)��pH��m8J2�'���4���Y�E��k�!��e<c�����<�������n���v�~��Px܎U�/�<;==�P���l
�K�Z��ӹ��y�b�[N�?�,ʄ&�x�-��7`n�)�p��GDZb�9o%%_a�S���E
���^�8"N���c���B�@�&'[7�w��������>�+-��"^vwov�[�U�W���	��5\��;t�;��qĉ��M�~ُ�ǷC�O��0��g׊mB�i�h���C�;���6MM� N�[�Ըݒ��ȏZĻ���=���_��w��y�_>��W�����������_�<��O/|��M@
�?]�у�?ef��X�d�I��<7���)>ۗ�bW[���S+xqq]�Ě�G�݅�n���;����+�p(��|��~��n(���Xc}vԨ���G��j�-��(S]ٓ���^�_�Sw�Xe��ʐ���D�����>��p���C(v!��v��u}a������y�y|�1��3_��d�4]ԁ�*��MR�z-
(�!������aͤ���|�s�J���kiL���kj��3�b������;�ۼ���d���.�ϳ��B��	��LF����'��������5n2�Ɯ!�('�����|��K9��$���*z{������Í���g\�*���`����Y�=�g���0�������<��c����RCo��^��*g�Re��x��1��ښ���T�m���v��Ϯ��!�v���+��m��";��Ū=c,�<�����^�>�\{����Na����E����!�t�،\���R&���꟪�_��)�����խ�����VuXD$k�N�	���]b�չ�����H�@�����lIؕ6��z����D��2�&��R�c mo�>�S0[i����F
=��d�T��{m�	];x	f?{�r6Y�U`b�c e����#y�mZ�}��#�W�4���C�8*R�0��O�]�����]tE�����GB�'�#�:0�����Kg��i������W���Qq�z���	F�
r:�G� vzn��/��������T��]�@Q������؋ͰR��_f�2u�vQ�j5p瀙�Aߪ�í�n��6��I��������5"#fg��I��Ք6����0��vp����ў�y�@�fg�����Az���	̌p�����{��#?q)�|')YiS�m�)�g'�\
��d��n�?���\�Vp�"��N+K�p��#Qŉ�(L䘉z��n�S�9��&B��>}��L���A���Nn�M�n��e����=;�_ZN/~�G�����(���݇jӦ���5.��4��s}�ayN��h�2�4�n�c�(����i���t3Z{��x�4%r����Ue�p�ODh9 ����Ay��nz��oS1?
�
���اcwH��=@7܃�U�_F�����苭 q��}Ḟ�(����OD�Ri�)�U�!v�]L2��3ݾ��T�_���\���&5��ֹ<M����o�B���J|ʿ�nJ�b�64��i���Ӈmv���?�ʦ52S�PւG�o� �ãx#OO쇩�m0��
G��e:��~�$=��%���8c�Q�[�w���v�Jr�9"Ā}���!��Q��P�%C�jl-4#v<\�*a��ӉГ�C�y5;�\A;����[�6�B)�P���2�%}v5K.�ű�{!���C���CǶ܅!$!��[���f$~cHd!��b(F��:5��y���g��)����%	t��:^l���� �o8gx[NԀG ��!�~��)�_����QP�?>�:����3�̭�6] S�F�Mg��U�x�E�d/��ch~�b�v-�ܧ�#�מ����CL�0���]^�T%���u:�ȀY�|�:/��5ۀC��O�~�6��N	�©�ͻ���y�������Ԫ��<��[���Z���?C�e8��F��+1���7���=?�q"c@�	W$E�&	�f.��Kc_�����̣PV�Sn���ǵbS<mG��,��g�ԗG���ELԠ�M�s������jX���J[]��ǻ��-�v}k˽�W4���ٵ�`�L��x����*�z�ST8����������/K�)���?�����h{ Ĕ�ݟz�u}�-���T�"�9O��-��F�,����_~����R>9"tj|&^��6�\h<)h���Ji��!���x~����{["zzh"⃺9S�vs^��������8s�wɢ�qy>���Q���?l�w��]�q���/�c�2��e���z;Ź�𩮶���.G���?PHwȘ������}��[���=��3����c�
0�$Zf3z�RÕ�i�ŴQ�O���I�W�4�K��b��-�����8ɶ�|��>�E�՛u�;��&���T����@��A��L���z���m���?��<#����ҡ�9VD�( ��������@��c��q�і�G$sר��(������?�䌕��e����!�Lˉ#��L����h����;r�3�t-J����p���6����6�
�ח�2�NR�}.f��u|O]��)���bɰ��Rtf���TX�WCB=:�F�eA�zw���:~���Z�6�����$�7/l冭7�<ǌ(��Mc���3J��5J��;��0��p�W��.Y�N�%��c1$Y�`����H0wD5���� �|�>�{,�s�[3���νK	�u2����3��sE�kx�1���xJ��`=݃�Y�����yXAX�'�'��LdU=��G>��:ܿ��x�r���v���Y]$|N1]ק���H���"D�T�s�z�C�l��B6��M�D��X�oΨ�ͦm�-)w�!:��:v�1@m4�$���&�v����Su�t���8VEn��pHe G�5���m*�)�Np��_����Ie�/��J�� ʇԥ{�z%�ֵrd�
����� ���fH\��e���g�D<m�;���`Rv�a��e��"I�a���lދ�|7���*�,r��	��)&V�\?�(w�u'�;(��ʶE;�`0Vj��%2��R���??{B�e,�j`�D�� f�O�;$+O��عvL����/ԅ�^��
�ۍ�gO�L������h�\�W��������	��]wX:U;MF�tJW;;W�
�He�6����n�f"a̋��\�2�4O�gO�&���a�a�FZ��H�J���wCO����/�,I��#�:p���ԏſc�,���hz����[���?����� ��}v�9���̥S�O����M��#�
���PLe;d���g,� ZRiWU49ܓXI 7	��O_��?�~Mr搡���10�/��O(�� x	�U����k�u<�!q�+��0�x�<Kg-)i��A� PT�����k'�[�:�Iܐ�O!������rBw6y�~�����Խ0�����8���(KXm��9V�b(w@v��qO�]���4R��?5�����ޟ.� �n�o��S�?=}g��h5�E%*A˃AO���g�Z8��v��` ��I�J���Q�y�5={�6��= |1��B�6���rh�M$�#�bj�wq&��-�^�R����4D���/&^�}��N�F�N�]1J�V���0����/����AɌ���4�q���S���\���#�xǰho'yV��Z�|�Ph�5��x�n�d�@�7�d�I.?�>�g��f�xȋ���[���6F��f~Q�ݎ�d$��r9a�5��#'�՜du���W�Yek�D�"�~�B"���q%Έ���j �j��ʢ�ͱ@�����l~7�/t���2�ǚ�)�|?+}{UX��'��,o��᡿EH�[�7�X8��=���|�Y�d!�t]F�;�Q�k�ʱ�x��y��|��~ĉ�Ϧ:+T��͵��I�*�$7*�[���<�LB �
!��Z��
����
��W^��
Զ�-�+�
�6������<�%I�45��UeT��	z�ol����ʨ����� {�?W��h��ICڊ����h��/����&�~�o'x8��H�U�Ƶ cˍG�7x�2�c{�}#dV�\��{�o���h~���bq%�h���h4�hb��<���b�����=�z�jnt��N�]��7�IɯQ��,�_�U7 Zt�I.t���C�3���o��̑�ܭ�ڏ�t!�i��$#1W֯X1�nCl�d�|_�<�%�}Ɩ�V`c�\KK���閯��͉�[	hq�;w1AI�ʮkXqӏ���CΝ�	�+"��s���'#�>o�����������f݇D&$e��}�ӿ�]��"+��r�{���/VI�:)���Ã`��@M���!2�˟]����k�ґ�����Џ����������91�\�_�P}%U��(T��s�죺mi{��'8"b1�A����͚���g���U�b��l#��RBbO�.��n�TX��E�=�"�k�D4oc�?y�f�����ƃV�'�}�-��=1C�4��%�)ݕ �2��l�oa��yh�wi䊬p ��bY)�����A���/�Oy��P?�i:V=��3*��R< ���"�c���.zKr�L]��/�wAW�xupK�B8�W4uz|�����<�o.�������'?
5�}I�y}n:�̮��+>w���qE8 ���#�������b��g_�8�з��!��C�ĚQ�}��Ԋ�]�"q ⋘�1w`Ѫ�9 L�0���{/r�� g����H�6�a
usj���;ޯ�/��r �ϩ�mH�БL��z :���[�B�>������`��YU�E��5D�pt���4�˻,��=;���S#׬�G�$o�r�ty�f�1uy�j�dD��<�.���_kr�ƹ:�H�,QH6 �bN�x8p�`�۰ڒ��[7�[�N�w;d�o��tB��%�,�b0���Ю$�/֤Դ����8���:o[��/�R��z�|t[���/�k������[�]ˈHd�ɌYp��؎�O@k��o�z���c�n~H�hE�\Y��8��6�2� #N\&#�u0X�˚���d><�8�⫄�7Ѯ
x�tF���W�a噕�)�Gx�w����v��$��Լ�
��a�¹��6��۽�`_�du��%%�.�Q�BM�A�"lçXx;b ����U��fф�B����ZD�R��+���{~3��#���D�����(�ފ	������Ú�c�,���*�ӱӠm�B'��wr)����o'W�%��G�}>�"ڋ	��V�4�w2��a�T����DO[>S��sd��������7�m�����t�d�+II�,3��IIi�3�rU�t��pƞ7~���m��^�t�%W�4!j<Ke�����h���.���A���y�L_�\��!L�ҝC}��/&ׅ	U�MZ��F{�p%�[MKX>;m�d��������,f���>��,V�<d-��5}�Iǝ`�.�-	�7;�S����F�+����K�cX��8�O� )����~��!����V�9�Qw�����x�m�M��V��Ӆ����+��8}5���/�hF�
�U�fe�JF;�|�.4��Bᴱm��N��X���r����:͠d��S�*���e�ET����_T%�ǋ�>ϫ�gެL,�$����X�)p �9�.D�2˟��N�vb���|��!��:��F'��! �mK�6�y1�2e�.�Ƕ6��3�u%�p�6k��eȄ4zlH�h� �9)�E�oX�`���7q���|l� �,π�%��ʓ�:��z^G������ʖ�L���Ήk�*Vy�#��Nʒp��?����T1�ZoY�e�Z*�s�eHF���/�'��
�\`��G�;����kI_�F�Wo��S�,*��;5;�j.f��K�F�(���n27��Q�H�P�9��)�������Sa�.��Y<vy�m�Z!�>?Ɏ����'c�^pќ�oA��l�����m�F�u��&�V/{b��)��E�"�� �G��':�����*�壈�+1F���O������'�;��[��9D�������d�>,�l���u�I�x��U�p�/��H��o�uH�h�5��E{W�u�yhA�m��n.k���;��~��]?& ��?���:I<2mNE)��M1J+&�����[���_�,��$J����C�ܞ�jqb}��|�<{��nT�;|Ew��J�n���bF�x��>�K��6cI6sq�7���UϾ���G`C�&���Vّ������)�������r��1ӿ����Д�JBl����9�W3ɪ��n򤭔�'|Z���� ���:�7���	���}	�f�]�����E��OZʣmGr��#�c,��o��J������*��eZ-��ׇ�1Ra���:�r�����i�=q�\�3.�����C����7?�ӧ�j=u�:6�<����W�}:���:�e\����H��?�!]�
P� Տ�C����b8skm�Lϫ�~�ֲj`���o�!̌����֡���<&�{����9U����'�� ���)��ˊ7�;�Qt���!kP_��,~�T.�����tAb�*Q�z�mŴ�g��� 	%�a�� �f#��r�T�z(8�1>.z㡹-xh�Tީ�
�:�
�T� �@����(d:�����Z�#���l��>S��h)z���h�C[g��ٿ���f*�Mr���Iu��|ɋ�QA�o_�����}oo�\7��ʋ�I�j6��/�����ȑ���,nY[^�鑳f�I�A�>˨w�=Ki�v��/dwn7��[+m,�c��756�he3&�>�۞��S��w2��'������V蓋�n���,��/�Х��BzP,A�ԟ���f�-���O&4	i�Ro>L���
P��9���d�;+��hџ��y߷���	W�}~&��I���y߆���Ͱ�[���Y][0	�^*�:�Y�D�J:�o��~U�:EZڂl�LC]Sc�](2.���XJ�s�!G�d�a��s�ł�ݕ��o���s�U&Stl����s\�ژeA�\�ќ���Cu�K��y�/�r���*��f�sdO�~�=^c�������E���u�o�]^�4�B���E/��+k�V��(A,-� ��p�mPڜ��)DI솵�z�sl���f+��~�M8ߌ��Y����2�αۡK!��>�#x$lv2� ��Q��&����:�`�2����g��A�!Y7�zP�zJ�CFj+��?\����.o|��w�
<�$Zr��9!��o'��[��9Mx�{ˡ�z���}Ȍ��a���q����b%�$���^�i=��~5C[ٛ[q<�[�b��Ɉ�W�6̇2�\�&��¼���G�ix�W�/�/i�8�n4<�ه����{���dj�
�ș���2�>nw� �3��:/Ԩv-:P}w�+�v�{X[��-![��^�uH�b������^q�&'k�ZsE��N�{�W{�Ez�sb����m+�۶�3�0w�u\y��aA�}����˫�I֩��Z��� ^�w���n��*�������wvv��[�WC<�����VS'��"#�'�v�5���&;�ة��eݱ͈7����~���j� :lJ^p8�D񽽵aS�s�Ҕ�*;��邴��Y���xl�����Sm���7��S���9S��,�KW�c.㳎�H��~w-G{g��Y������)���?���7EE%-5_�D<����F�v�W����m6W�Z�L�K<�D�ȝ$�94;��*%�S��:+���r6R��KP�h��1Y��i�:�Rypl��~3�|w��|	�q��Qw_���k���h�I/�E��	�PZYX��N�as�El�ȥ�J� ,d���ɸtՁr��U�����=f�%�gN�����^���a�-`�NZo��$���'�jJ�@>Y79����f���T׼@����AL�Ё�\����_��~��蔎�7��ݓ�]}g�.�V�����6�E��8T��50�hb����ѩք÷�0)8]]����T���[�g��k\����~b#�1��R�>U���8�U!�������v�ȓ6�'�v�Jy�	<�/4umyڢ���e!=�ǕZ���s6ǆ����&��՟�����w�����x���ĵ��1qO����~���Mيn�Y�8k�П���LMQ��z�?����}�M��UHʾ��D/�~L �s��{hTbl+�s��w�ߐi�8�ח��҇*�AF�m��9}���_ϥ�ER��k?���::����C��Ԃ)���_��8��*�P�@[}M���}��>d��B+t(x[���$k��{���R�΀��X��o%��odC��&����Z	��ҁDf�r�r��� .���\�FW�r��*NJ�E��|R&�UG���<��=nV���o�߭om���i��U3vV	Z&]ual0��;՛;�(b?��z6|���N&�vtn�Xgb>�3�_�6Ш�So���s���7�7�m�f��ı�Rah)�h�#@I��;��}��zqԅ�����ͱ��¾��/��0�ܟ�LR���e�����a��k��à�"�Ъ�
!�n�÷�nd~*��6�u>30�C���I����@���zv�\����%)�0�؜��\�O����u&��r�~_�� z3�������jy���,�"�+�P!�{yq#(�K������YS;Z������(Y�*ī����ri�)l����o�DnR��n��kk�f����o>�l.n�_��5 �_��ɽaT�Ep��_��>��2�������R�(��Waa7��"&bː�����v�(�ߛ;��Ǧ����(�rٓ�������s���QM��s�Ks^�Fxg��'�^�x�YE��Ao�X��0z�RM�$���u�X\Q�����-�n���H�&ܣRx%���/�h84��mZ�^�WX�'F�Ҷ�n�s���
{���jv�|M�0)mg'Ȉ���r}k���8�&�w�;5K,*�d�%Ħ9J� 9�ʍ� '�d�T�(��`��C]�)��Vm3g��Y�rS���ٷ����h���l������Z�#v,..�>a��R}h$U���s�M��o��F���l�����L;�w`�3���AZR�ͻgڟ�7צ�5;��?l���4���v��	�^�n!+##s�H��AQ���fre��C�WT�d<�p �V�p�L��%dԶ��"dՂ�ق��z�>J>hY
�����`�z�O����y&�щ������2V��ױ�L���$�+b���f���F�Vq�d��S�]u���m��*��^�"�^���yQf����@�a���\==P崽ok_���9p�C��_i���;`-����'�|�O�/�ai�j-���%i�g� �O� Z�b7�HNdޡ,�W�bn�	_�:���7\0I����(>�W(��<�����[�W�J>���>qӄ��|�:8����e���j���j��ʁ��mp��~=����G�&|�������� ����#}]� :2\8�B@k*?Ew�{ ����b���o�T{���?thZ~QV����M��z��aL���o�(�1ƽa�h]R;^UF\��X"ͤq���l8�ǣ}�S�f�g��	9��sr����_��4*"-���1a5m�kˈ�|Z�)��W�"�3�˲�]����cG���b gƁ�fgm:�=���^�ٽ�h&���<�^]�Q��=,��7�:.T��-,��}5L��?� P#|�E�����I�rQ��da"��h�/&L��̯�̵�GP)���ϩ�cSNNiHX6M�[�eܵ`��s�.�"��a��[����ܫ`�q�N���e~���a�����J:�0������?7���A�,Uub *��òt��55%ǹaWH����>k��7*��~�|����r����z$���݁���JU�n,k��}���_��ȟ�%|#G]��P
�Ҥ1���:"�����U��h���u�	���� �5����k��%��]m w�vzQ�))ٌ���)P���ʎ=��Q����}8���R�w�����x�� ߪO�y$�cl�����¿�hp23�m������)���#�1w���4A�j�/��`��W�X-_	��[f���#���ƺ��������e�6��]^���0V��k��J���L����v����2�����ё8�n�\.w {z.{!�nc�#��tx�V믮����2[�⥫�(���X�k0VTJ�t�-���L��>_�C�<�n��4g�S�ձ]L�2hf���(��J5*�g�V��1h�X���!������O2$������Q���z���P�t0�a�O��V���;OO�n��*?����O%�e�~�
�!li[՘�� ���N}��*ez+���qѽ�Wfze��DmM�>��W��Wa[o�a�V�O����4�[��ɝi0�*;���T�
F���>�42F^i.�:>l�s�L��߻��Y�Z~/�y���_-�C�/�����.??,I�pO�IQX�h=g�_���=�;��\�w������q���J�}B�+uH.<%�j�G�C"��%���u�����[�H�Q0҃��=5����3$�%GE�eL��;?�3ߦ�ä#�����y:U}q$�w����w7�{���=g�"��1�(R]U7nr����d�,�_�]�X�y��U�џ�{�}����.��5f͎�j�9돲��BܯUc�(�Fi"�&_+�k7!��C�� wl�b��?!)UI�P�p(�{��P͊�̯���Ϭ�qk�� ��k�j��T6~����(���{�[�e]pIF����h����ʪ�>;��_ЈVEk$𮔖N\dx�C�0Z�L�\�2�#�N9~����e��v�����|�� '���J-'����C���'ζ�H��z����Mʩ����R12�w0 ���t{���M�VSw^&��l�[m쌛9���O*��05;[/hhp�Q������v �;��ƽ!k8�?��d��Yc Nm)si�<�S���5޷9�4�o'����̠��������z��j}P�7-�X�#:5�_b9�̬0<�P�؊�oip����_�q�"��b����6����P�ʪ�G#��Yu���$�.�Je����d��B]ZVB;��Wm^��iitn�]CW�U#;�l���ϟ��]���"/FF�h�cS�Z*���������!I�I������Uw�*4W�E��8cf4���K�Ág���5lF��P���;pQ��=C�D�!+��쌊���x�޾]QEq^SAHt		sɧ�lC��[^;&�J,<��j�ƗNg@Іv�_�s{��o�)��)�W��|?F�o�k�g�V���-`l�$'O�k�F�󆲇.��x�yE�O�vz6��5u����g�<j��y��y�,K=��J*L�R���4#Z������n녻j=Z���G���G�*�ƞv��b3rIv�M4-� �Q�TL"��Z�1�	���J��5_L��q���ۺ���<� O(�u}x[63�*��Ʀ��Y��ũ���E��'BR�,%U���͘������j�Q�o_k\�Km����de���%6�r{�3�R�B6��Z�
;�ו����j�����zX�S���L��(t�\7��C����	��_p�Ɔ{`�S��}���p�X�?�eKz����`,���#uhk�^�x���T���w�h�0�;���.�<��%vW�p]-�ʺ�%�������$�s�tIO�F���=�� �ǎ��߈�5�h�65�]�gS��5ҍ�c~R^� o0���#^_V|\8����Ԙ,L�*d 
F�A���.�˻��Y��@A�3@e{�@m���Xa�c
h&D��(�7wgu]�^"�i�pe�����s����#1�L��d!�ѳ!ݎ����o�O�~}؇�;lmĳ��엳)�m+��ᄮ�֤��c��	F>ćb�Q�L�jR+��.�׆��+����%��z��u+>wD���	vқ�JH=� �4�<���4�_H�s��[^T��G�@��'������uovo�w$L�o̢ퟫ���".�,�~@ƫ'����fT���0s���x��cr��a=&����I�������9�ʂ���S�9D��}�z�h�2�pѼ�GDS��]>��^�l�j}
z#F��<���1���������e�����v�/������#�G�5ݬ#��w5�_P$|����;]/��d����ag~�[L]��gi�ꦽ��rA芧�B_��p�b�;7b��%*���F�<�η8vw6�K�Gg���f,�_�|s8�׼��8Γ�\W� �z���ܝ��)&���go��gD���xq/�ur\��9Us����cԠ�^<�Ը����`�F$e$��W�V�:�-I8���4�;�|'c���LȜ&�8�e����0�'O�O�}�*1G�B��ںe���7��b�ު��v���"8��}F�[޴�o7 _�������Sa����u�r�[���Y*D�b\p�x���@�h�ÌÐ�����-��	V�a$�Q��Gڕ��}�هQ ����Op�K��T3I��e��a�p�~���~��nfػP��V����z�j�0~�9��x>�C:�N#~J�W��f����֙Uټ�6�̛;u�����I���sX�+)}d�������2�x�`oٽ�=�d0���Kp�L^�ޙP~k��U[�U��>�P׮u���(������)��B�A�˷����t����{�$�d&�mM �
���1�lZ)����v�G�~Q���Km�k�|�������A�߽-��'Ev�y��3.��m�c|M"���c�g�����&��Hޠ W3��"��qk����@g	��5���cx����D�(]��]�������c�t����:ⷺ��'��gX咩�߫��\����������X������'���=��E0���O6'���'l��}D���o�,��vEp.�?�:��`$2�.�BԺ��f����	2|k.����Ɣ�~��n���Ѥn��\�,_���Tk��MLgǪk��T�n�֜�j��oF���!a�A���m3xz�G��>	�Dүg��vwxIB�w~��F�����^7��1��>
��K��f�~M���v>��[�*/N��$����37�3$�\y�ơ��s
q6����bFzƉ*��_��!g����j~2Z ��>�>�KɍF^0@�`LR�S�������'��i�=����*�ن�E��2ƺi`�1Bw'�WӨ1��j���[��q��	���]�C������	wwww<8�����>�<���������k�^�z_�ii:�Ɩ�7,z�m6��%����6�
��SW+>wOWp߃K�p��ǉ{�S8跘����{�M���~m����f��*(���/��3Dwp=ay������-���cJj^K�;��ǧ}�3y���͒t��Kja�����K��t�����3}]ۈ���5к�D���@[ֆk�;m�h&�b�7;�\��ɗ�rP�׈�,���w�����6Ӛ�	[7_���7�k��UAn�N�\�����1�)Ⱥp�Dݎ=��F~���ƣ��+~S�ư�1Uw!��/��#|1~OLvk�6�/��?b�v�e�Eك����o~h��8@��Bϕ�aly��p�`�.�t�#W�vn�9��;�y����ťm��R+��+���vm!.�����b4���'�_?��X�Kw�FTsD��{���
�hqJ�,K#6'�>d�}�k��!=tzr-�������!�=AzҀԔ�`lˏ��N�z��L��'>ǋG�_�5�܆gj�����ŗwK�uWO��>E]�A|��!�����(�)��ɰv���k9�F�7��;ao��ךA�Nt��9K~���}����"i3>!����T��7��A� �z�؇y|��1*	�bʩʲMyfʷ}��.����|�c��
EV�����A5�+�4�sx��ݕ/pͫ��l͟84 ��M-8
YSa{rR�������C���P�[�8!�/`�>yH�q��ݠ�B2���.ō(�9I��[��}�n5���ά��:O7nSrO��0^��1D������ ��-��:6�������Y��s�	�����i]�e�!���e��o���#a"
��KF\�r���\�xx�\5= ��/v�O__����ճ�fO{�N�^�bF�QXhQ�@��}���햐�>�@'�@/탿�7��U-Rbh#3}K�7��	$g�(QX�Mn1Oݟ��h�踇C���HV�F��cYICzW�Dp�%�ѷ��&Lg�;S,�R��E��'�r����>^n��l��:��h�F�;!8�5i8C(2_��'&-���-��Vw�Iw6�v}��	���M|R!�Ӷ*x��%;�5կ	<����^��5QR@�D���wq�R�i#dm�5'��!��X~	FJ�0f�Cki�����lq<q�W!i��ڊ��w�t��a�}�i�9��PY���c�95 [��h,h�l�k�Bzn	��;֨�.LZ'�<�o��R&�Wf\g&�0Ɛ-�(���5��5�\�����#XGW �CF��W���E���V��P�mC����?�?y�D��l�)�~����0�6Nӟ]������S�����XiA������l?^%d�� ���ݤ"����o{Ψ��l4g�1* 5!�]z���Ǔ�1�G	���W^�6,�&���W��?(�����)��8�
�&��D��8	X����k��7>H\,�����)�PЁ5��+�eek6�`׵��  ����g�#�	��o6b!��xL�(�(��H+�}�����Ґ�9�D?�)��44@���]Y�ꐪ���7����^h�&;\�+&\���4+�����~����w��d�.���9�U�}��� |�D���%��<I�-���j2Z(��=�I� \(�-��ĕ��O$�+����VZ=�Ḷg'�Q�������[>R6��YZ��a%�)%'�9�,�Z/�Y�J��6��8��$�Lb���4�bZ��@�9���hWRR�(ط��2��C���ڱ������ �O���y��`� ��2� ��-٠mgĊ�`y�EWhO�A��pn|���Y���Ӣ8�#ح�vd(�Ic�@�Wx��A�x�T�79j��^��PV�%5��̟��a�S�"����G�х��hH7̉~�;�N �i������A5�J-(����l(A^���Ƀ����'����'TN��u�<�oL���>F �R{Y�~q�D���<�A�p��0�)"����#�aY��A#He��a�Ȅ. �ѰoW���e�o��I0~P#�R�}�vF���z���n����=��@�{Y�?#�PS�StLm� �f{�, �V���M��������ٜ��r��a�i�a'p�q$P{V0�x\��|�C�	��f?H�A�]� ���U�}"v��9uTw��M�R���ݏ
z뱐}�>�.��2���R�X��o\;�1Z������;�9�w>�^]�+[��8V���nm��)�MPd8*��ng���c�4����Mm�aK��n��Y��һ�d��#^<1�����4���H���w?�>J�V��t2���H���xP�?�>��_ɿ�$eB��������&�q![�w.3)�{y�e����':�x�F���@fc�ęj� �ab�\�c��-�V�c�og�ݝ�q�����k}Lb]Z����T�H����L���:u��;vk_�#�$K��򜸋��E�)ᾪ�ia#�E8=ľGU�ת���'�z�e1ö{s���1-]�����V8����^�T����!+�`tm�$.6�5;-�`�h<y{]Y���h/����&��<��4��S���r��Y|���fr���rf�jxHu���~�2fn(��)��2��79�s�nI�5S$�/F'¦ݝE���g��5�nN���cM˹�� ���\p�����i��`{���L&�u��5N�1�p'����\�;w�\E�uL8�w  ��xJ����}'m�|?}v��m6b����$��MR��?ʇn5�r�t>_4�?�����V��Xp�׵m"i�քnU�Xh�nh	�Y�G�ո^!�#���[�2 #�C�S+*]ۑ*Y���~d<]��R��#�Q1)���ɷ�n5�ר�n��wXm��\�R����bv�ŉ�˂����a���7�Ǭ�OgL�T3�Q��A,��6��t.�Lh���̹D�|iy�m�#B��B�@Q`������Їuo��0�=}�"D�<Z���!��y4h��%��c �Q�D`���[TN���8z�,=1���:6v}�S;�e��l�^��P��2y:��Y����E�'��I��	�*0C;�9Wx�d���$�%ćv<Fr�e���D.ݎ���p���b�����5�2�s�-������L�X\r�X�7P�DN��,؏&���H�j��U�N��~����S{竻|�}��I�"�VP� (|�6�3q�)�9���J�FdL���%{-�.�_��.yo:�	���ŧT�Sqm��í`�e���bͳ��y��Y�f�D�E �9�o��>�1Tn��g������?���i>� ~ċ��p+��
��� #Eiu�6m��q�k�rV2Jzˑ�����h�X��j93��!���	�N��8�w�Y�rC#W����N�A;)��a��.~��Ɗ�i��߳�ʤ�$c_��C�
_����3����z�~I�kZm;��.��m���eeg<)�>ړ3m)1��b��xQ���c��pK��XG�q�A��ީfflB➎�s|V�įP�����9c��e�o2��B����b�n��F�a��歩x/�vC�R�����{�;rf/��D���}	2�9�ۣ�����ϡs���|
q?ޝ5=?B����/�S�a|��@�Z98��]�u��yG�wk�{1)Ǫ�O°������@����g��H�_�scڭ��Z��e��Ը��r�#�,��������	�u�b����MN�T�䆮3��d���#5ԓ+ά�^/��� ��bN�V�q�z��pK�kzx�}����B�6g��Ev6S��7W�A�4z�"��Ǡ�ыj�@kA�K*���w6��g�����$���Ym�B_�O����H���l���g����ΣU�Ņ��cדV�w�8����9]
:-Fܡ��w��+�)�D��������co���̬���%��'ge��D���QG��+䈫��;<����"�N��n?���6�m/��&�%�BIB�Il~���+��^ l��'Z����\����J�ɛ`�'�t~F'&\Ho��3�H�n��	2Ȩ]�.��zr�|��|ޣ2�K����,���������@1����Y�)��i�l��h֧��ee^&�HF��EYM���¯UEF��̒�w3,��5%�:�I.	B
{�<s%���b###��0q�o���^���>��:Ɨ�}��6ڝ7�J�>dn��~�Uk*�~3��16��/d|�%&l>��@Ѝs���K]��ٵf��1��L�:����{�?�|����F�/5@�"��S�3z˛eV�����Td~R�������ޛ��l�N\���Ԋ7����jJ����l�܇�,�7N�������(�/�V��_��<A=��(��99T������Q25����-���uH�P���7z.e�7h��٬/��踙��_��c���]W˗jV2��&��,ۺ�1SUl�H�9z2eݓ��U/?���R�٤��cr�wPs�ď�ĘN5\���������2K�޲�$4Ә��e6l��T�П�cc7y�-̕.���e��;�f2�NmB#^	�?ؒ�t�H�%���in�VFo�����V=̵iP�Q�G��~��;G��g�II����xzҹ@��<�40G�s�@r�Θ� Ѱ���4��6vR��<sG��v�6�o����vJ-�,jѲ=)fcߍ���>]��rp.�l���:ٻn��(�A�y��-w���\�����L�{�����J��GS��
�H$�����G��e�;Q���VC6�����CoXD�wG�R�F��F�̗D�|��t����Y-�>خou�V�u����[����/��D�#bbm�f�P�P �V1w-������V���H1u55X���%G�3�u����E��W_��V���U�wY��k��1��7����c�?��l�.�6$��=�q?64���S)1[Rݝ�(��<
 ܑ ��,X�����D�y!���w��ϥ����Yoyf��7��|^=x]�zfz����?�ߚ�5��@���p��=^�g�{��SV�qWn|3��c|0r��}9)�҆\�ߑL�x�@�A'�a���좮���&�_66�XO���ǒ���T���Y���?�Ya��F�T�����:� n��A����R�EABv�oXG�])Pz��l���J�����C����Ң�"tl-�=�?hq�`�'%�\9���7��w�P ��q1�t�ɗ�1�8���i�l��jB3�i�G���z�"A���\������+����쯭~8[�{�!�K�9@�������}mTV��z�󣗛vfj�K�QPQ��N0|�4��֜�L4{��?�
�|q���w��o ��%J�F�a�e��9K��ߣ���[۟��B����Q!�#�W���t����S�-���������|�|�IBBv���jD���A�r> al,&��Ù���O��=�ax�-
ض�X�w�$T)�.�񑊟18�:}pry�rάB�;����"1g~�/��~��ь�����+�ҡ�d.[�z�}!z�;�yJr����ˑe�+Ypzj�&�2�#�=MS��L8�g�ȯX��eYC�*w���e����-�>��z�9Y���ZÕ�ſ��>���Ǵ�H\����NWW<�W��%�s5,o�[�}hY���5�{�Z�&�a��yV�n��E��>�~�<��$���S\*E����8��2o׽����V����M=����]@sC�6��A�����Ը����F7J�ף����Ν��-��r��i㭕���T��.dg���O�e�m4	ֺ�@��L;^;B�m��w���<�����1
���_�����\Q\���S+�
�|<!�	�������i�E�D3�3ي�݅���O��G��.��?������(�vI�/8��C,��
$ �������.�/mm�=Ń�:�]~II�~+��2����fr��U	�X�ax��e*����L��Xx��B�/|���O����a��^�ϕ�����Xq���ɒV���=��n��@���m-��T�?5�(�����*N�][i��u��Mǝ�K��u=8��x����JM�&Z�iR̕�l,lo�堚����u�(�;���)�0�P����5Q�"�
��zlj����o��y{ߥc�#�W��ݿHM�����n&���a��h��K�`-3�￸-��x0I�?q��{�|ŀ�&��cV/ݖԌ����xR�AX/�ՓV�v뼩�����z2�����ǎRC�F�N��ȟbB�:��U?�F��p/䨕�S�2q�ɭ'S҇o�ګ/��"Q���b��|	\j��3ꛧ��^K����!�Vw�?����x_Y�����2��<���l�(���Y���g1Tv������u���+�j]���hPL�L�>��T��Jz�!�ޔt��҄�ţQ�m
2ǂ*��D&X�5���.Y��������z����z�>}S9�9�ۉ����ݘ��:���f���A����#j2P��:�9x�~�|d��e���d��A��1�խ<5;<N�lPҿ(��vv�PIZ�IKF���P���^��kMHӡ˨QwR��O�sL闢O�?�ĩ:�/�R��������=�6����ȉ�����N6 ޻�\y�Z=�&���K�Z���Q��O}0��Fƃ��|{�!"W6�Py�>M�����@��ۉ�{E�1�`@��@<ot�ڀ�s��4���*��+l-��AH�Bv9�����8�Ҫ�О�c�"B66�&��٭e\����������(�N!�nZy�]�!�dU����~�G����ц�d�!�.�� '��-��u�:���{t����߻:Ͱ���P�j���S��dB&�������(X���J\F=�ޘ�������K���i��h��择�Bq�~(Az�9�_&X�F��Gn��$d� e���J��5�	�{��2zm<fc��&uD�{q�8�@���,��⚰��� ��[[��$��#x���̉8�E�H�3�k�}ufP9L1��6*�a�0���[�C۵Dq��,Z��L�A���
���e�#���:S�kاL�z�9q��K]��V7u�J�Ny�1�z�7Tw�+q7}��;��'�ϰ�~�^8�����"��E���!�e7Bs�/r�K�h��5P0����P�����w�|b{΢����s{�D���l����M�rt�-S�ҋ�w1������
A���g:�5��3 _�š�
-g:���9�W��
.*$�A�`y7������0�\
�X��_ z^�8|3<���J�B�#Ȼ�������]�H�(`ױ����lȿj���MBӠhU"7'4���
@�eP5�L8�Ӧ3��L���~��c*)R��[��R���5�'���0�}WN�݆�H���6#V��,�&��������ڸ�{}RF1f��NށFV��.O��Z;���i��-7i��?�o�p}���"���Y�ޭ�BwI;DE(�+,�(�dw�:%N��Vf�X����*vqRE�[e��N� �R_�Zܻ�'|�4F�~^����CJ���L� ��s���Ǿ�S6���l��� ���E�D|
B3�"c��&*��++%\o���a� T"Բ���"j�"���C���I����Žm�ԍ��W�DU���w�O��h�����%���{�{�)-/_�[~#���Zx����d(��~~F�����T���%�!G4�1�?�;z�N�<�q��k����\�U��9����3��N�`mvM�w�o�3��L����8��rx�ڳ�g�ߟ+�_k��F��^ �;�&��$�=���Z��c�D�B*���gs��c���8c��XskȲR���5����a�>��-�)*f��LOͿ 6��2w>�'ٽg&����ۃ9�/�@l#
Ŕ�dԽ�(����K{Xb�u4��Fu&�[��]�,�m��K�G�(��uwE[��Y'ej{/�<T��Uϥ=B�I6M;��:���y�o"���;���\-5�2l�����xX�;�R���u8�SW	�r�� �/��>��m$z�Ow��v����Ƥ����Y�l�)�~����g2���1�Wz̸�����<�g2:dU��9��)"��.��6�k=#}��E�b �:zqo f�w������*�7a¢�>����{02��^2��iL�r<��E����]ꇳ�F�H�{�x�Z��>�{n�q�����'�Y{S�)�;�t��0ĝ��V��p�y�[ٛ��ۘ�@a��Gz9�&[�{R.���e���Aʫ�����Ts�x�:O=,	��^�!
gw��w�i����DL��W�Thwx��{�due!,�,�zڡ��3`܄��u"�=/�>�C_�}��ٵ�%�rp��u�L�Q,Fke�vl�"SD	���UMKpϴ��d�ko�KD�n%}h��w�T�8���ni��+�Q�}��ʙ|�K	��7�����C �=�h��|j秩J���V�A�	|������s�P�+��l�"�rd�{{�Ӛ0#�2�ȌY�-3m�L�um$i��M���{�����p�)��I�3�H3l�(}����{F�_UxE݈�qPf�iT�E��&Ô�ST�>��OFC��'�1舘�'��h��r����z�;��?t�XV�^^�o�%7l��K@��Fg��f�=�.�<h�U��EzI�R����巈�E�E'����i\qd{�j�#������[~��Pq3���G�,�ˌX�Ld�ԝ��]��ڳXq R�)�.7�������n�5�*�!���Wߢ;Ez�����Y���7�ʴC?���D���	�W*��G<��ca�_�C�i_}"�tz�(|·�&�b�=��`ێC�Fi�Tw�X�ק�"_0f�[�V�moL�?�Oh�f��iv=��5��Z�
\n�-ŝO&��3�M������crL9�9�\�>t��Z�:|��W+�mbf>�Z��7�h<U����9���F^.0�h�����&� �$���X���V2˕��OR_�HT"��D���w�����qQ&%]�4��.n�p��梿�l����?0~��'�]�I�,��-�Iv�v����w�ʎ��;B/n�Ͻ��MS���Y�J�:�ѻ�cq���=�璬��+>]*h�y�З|�Vc�K��Y�{**VG��<�J�E_��3��~7�w��22�撓�[�*Uͼ�Y��.h��
�[�u�wCc���r�+���Z7.��^�9;�Y:���Ρ`b7��AT���L��֎7eƲ�^Bc�O��2�_=e�̉��kX&4�v��W�Ӎ{�wG�����}C�����%z-�����#�C�����K�fΟ���}y����j�e�4n�/}7Q�ICk��Iֲ{�����wN[J���)��D����6��),�_`:�{�_�'7
����\ks�k�Ի݊h��P�A���}x&V�Q���Ж_:¬|�TIq�,������ܒ;�@�@�\�]]k6����N��:����&>��UwLt���0���{���e�o�.m'BR%���w�[P���ho����Zlw�[VW�9�a���O�ko=�L��n��ϙ˥W j��8��ߓ��:�/=�i�W2vj=W�,��[�%k���RH��"��B��v�E��
�l��
�<[������F^����cn&��y�.Y��;D'���1����(�ϼ|��^�!5�G��n*��V|�%�lKNl�4��oKuw��^��%��>"!g,�����xrF�x;�`Bne�:������
>y7:�p���yc����#�b��V��U=?Z5L;50����Gk
/ʠ׬��(d��k�������I��}��׿.1��3�)�k=� ?T���R~�i�E�C¦�+�`^̏h�H��q^^B������b,���e-���Q�O���nz7��b�N�+RB��M�������ۛ�f����H�Q���Sַ{��`!-���n�PF�y��RHmL~D��S�&;C�Kz|��z~�z�vc���������c��1�ӿ8��R
�;:�-!�S�q�#�� ��n}���,;�Y��.l|Ƭ�4>�d>��r��9�曥Y�L,r�c����'~��Ȉ2���:w���^x�ZYN��<(�QGQ)����,����C^1&<��w��P®U��1�aakG��Q�x���X�\+Y��g��8*n&iN�.N����Ɗ���R�ܸ��eoF\Dl�$�Nݦ)�	'�-���l�e������6P�d��ʡ���:�d��y�q~���c�[n��ړ�����N�c�+���4ܞ�Påz!�$C��M���/ܷ9I�M����s��G�Uv6���������︽퇆���/�o U����ĸ�s�J�����x�2��K^X�N��
fE/���7�}d��1S���c�.���$~Bzp�(��m�������h�6�C�wN�W֦�y��~��˪ ����l�YY��9�*�����F\����$��?!�q��m����v6.̻,\s��d������k!f;������.u� ���n�@CBR���5x���my���-���~n�&~ZM��n|u���PE@�:�5{-k���:n�9Q�i"�]-�e��de3`�V%:���ѭ�O��ޕ�U������p�o����V�tȸ�?҄l!���4�mq�|r�����Z5�P�y��iW�i}��)g�>lt��"q�T˓àa=<���Qwno����&�Tz�m�B�������,���0w� @������Q�S�=
��4oH��J91��N�)���˧!!d�;���J�NW;����q��>zeG��{�sQqDA��,��m���'@P�Uqn���5� ���b�h�&��mhe������[dY ����3�JF3�ۥg�[��r�+����r���q��[ [�w��/��U1q,�V1��/�'o�(�Z�¶oL%pxp�&�
�ΖG���5����+V��N�t���:mY��6��"TK���:U,<�Iw�����D�K�.^��1���=���X��vA#�[Jg��;9��׊�'6���"�����N-\��a���db#��U�8��A.m���Ga�!y��"Dp�k��n>~H.RK6\'�]���@Xg������k�]�6�,�P�2�^m���YP/u���K�z`�gu��_��N�������7Q�O.ӑ�ʍ���iq{V�;��v �r�fL4�;��L��c�6ސ����n_��Ĩ�ézvyµՍ_Ep�)4�wO=�t�#�}	��E����~��c}{�����5E'h���M_t��bg��T8E��};��*����M�$�ǖ*
C�e�0�@�,����B�b�+��uАN~+�P\pvbi��b�� h�S�5�+�T�oJ�T�r��^�1a]���6���W���&<������I�Nvh-3|�KW�'�;��Z�S[*r�z��J+����a��x�k�)����4*1�q���L����{��Q?���W���ג;���%���z����zx�c�N�0�~������1���8�ꗂ<��^gSHK�2yF4��*7�iz���Xŏ((��A^�MR*��dW�x��:'Q�S���`��B��説|�ç�{�m��s�������S��c��1�y,R��*q���~����G\.��P%��cn�ܪ��l����r9[�E�p3x�����:NU�S����,�]AA1���>���I����`�b�$���=f��"���j$FtL���1:�A0��N���G|(���_H�z�����CD�Txw�ǁ��E~��נ���sʌ��n�	����1@6U������2^u]�MA�� ���l�B�"co��fީ��0��2'�����&W������VN�-3�ϫ�*�z��EP�	s� ^-a*�ځ�Φ ���v*���	:��u 0�מ��A���]�=�a!��~Y�kPhr��G��5�5����p��m*k���(�H{��3�R{����S�#��Hő^��,7����$��U�v4�Y��B������ei���!+_��-�'����5[�{�x�����&�*�Y�����'�7�tvc���Ew��S���̮�)UKf��x���]��҃d��]�a���e!Йg7�3"0�Tm+�H��35i�ʒ#3�#.G�HPM����/���/�-� ��-@�"&���+G����ŨIp��-��$P�$ f����-��e�?[s�*3,���g�l�U�JDG-��7Ww��-���4`Ħg�jCQ`|���\�E}g�����8>3VC�w-����\����9~�"	o��Z���`�oIy�����^�7�n{�U4�|t9���]=�©k�Nfw�K,���kM?�30;���SvX���-��G�Y[䷐=�Y�OU��&:4-:6�lv��%��>��"�QW�'\�V�/*���2y�[���xQ3��Xu�{��ژ
� &�$�"�yD;�0N@s�p��x�T��b:��`��Y75�O��tk�;��nDz-�ZI`'}��P����	Lkn���\<�it�[P�d�ay>����G��Ba���~�?�D�JM���a43�`�9�Υ[��Kv������?l�ŵ�e�M!�)�6G ~�ѡ�ҿTMh��NO|g}S�(H��Z �.�������|3/Ҋfo�`>�Bd�V7H�w:��G�	�g��n~G�ޯ�Y�LmX��Jύl�F�i'��N0�7��ZbO[mEmN���-������z���e��痂��H~�:�L�xS՝=Pc���;��W ;.���a��H6&Ԗ��[��nm�ݡ�3�걦)ҥS=9��V;�Ѹ�����y\�;����2��Or��h'�R�$�sk.75ByY��<�
L;K_��فl���mtz�?�׷<F���NӴA�/��r������(��-��4�L�G��{ߺ���^�g`3s�0.�=U��Gz���E틾��a�t�+9K��������� 6>mG�R`q�t�!�������J���'�s�:'��|�T#G���0���+Q4��zQu�l���"�0��Xvh��=4߶cu�eq��\�BTV'�F׷v;J�aj�
�1\.����]?_�N�8¥،��Y=x�=^Q���ZN�r�#��t��ш�ɍ$N�<�Lo�Y���Eƙ���g�[��TtU���'�$丷�0�c��2�������/;����N����m^�+z���ǣ��8�8$/��\H�6DNy<d�O{�kO�I�L���̄���p�֣A�̘ݓ����Z���O9N �kKg���*-xR�ݝ~F
�m��p�_ ���B���@O�������i	@�<�>\���j�����(ؘ�%�g�Y�j���a;��W�/]CiȬ�Y)3ܷK�f�0NU�".�s*�Z�c&���6�a�<�8��L.D����G�UJ�<xhn�=��y`�o�QO>��%�U��6/fL�-]y ���Z^��fh�Y
7�2��^��h�����ʭ��?͍��X;�j�E�o~W_Ve�y³}�K8�|0��z~�ObV��p޼½��t�h"ŁB_�A��߹=<�|��a?uqMa�bui~p�#�1�Nv�����d��kB���2����]4f�7��� ״�p?M}Wu�`h�W�>����ek�e��[�
�1���N�rۯ���ۧ�ޏ�nة��i���^"�\��w>�՟u�p�պ�u�f���q��C`�o�<"b>&�Ä*�>�ۄ���r�i�����󓘛�䧽S�r]J���1�t���2����f(W]h�.�5O����Bv㉦u���K^�ɢ��w �!�,�ڰ9���������_è�y���T�{a��Z���m$�۵��=���]�*�4����lʹ���(���2�������Ee�)�uk�®�,�!$�7����۪t܎���d��l���^����Q�Ȕ��c��_ہ��1���/Ϭ@2�~�з_��:�-?���O��v��Ff�r����Ɍh`��ɬWx�����$�G.�_�3�J�������J8G?S&
��S4v]=(N%X�'��l� ���1D���2��UUW}��Ĝ��	���Ő�V�����pxIft?��uZfjPtU��3l��^���,�3�|[
3�s�����%$p����Dks��<�2�~	}�b���LȻ�5s�Ң�0���,#=u�Z�9D||�I��w�.��yPA�7��y]Y��S���5����� �xf�_�x���%����y\f�����s�]�^����j4��ew�r��݉o�;��
噧F��^qF��o� ��U�۔�٣g�>��,.[���by��9�2�_�Q����2X�/NNN��l�ay��j����ض�5�|KnN�|�\vK@ǃ65�Q�z��x��|�_��Y�>����?3AOй��L�����Nʠd�����	��^/�����T2�v*�qq�|߲�X��eAo��7���c3����l|	�.� ����99��̪i]Ʋ������2�2�H�=	��4"^τ8\&����e��,�QG�9t&̝o?v�;F3%�K�������s�:��U��żv��4���L頨�N@�	7W�����޸�:�����e�W[�s?0�|�����R�Y:��H�.�ٛ����߄���<I8A Q�q�۠u,I��0�!�	�X��ӝ4?����3NT�^�ݲ���\Qw>���H:��uf�-SLu����JH�-����D��[�h�70ȩ��P�a��Sܷ�ᬶm'��>װY_����-���y-��#��_�|������OU����C�&�&�:~��1���8 ?R��A��4�(K�ؓpx(b������mgO����(���	�W���;��+�b�#�!�SF�)�b>:Jm�c8N�ah�����Y146��l���K�O��A�^a�۰�V%������x�Rbg�?������5�)��@ޛ�<�{mI9>�"A~Dx�pJpo�Ԡ�J��_�W�Z��Vn]J}I���=�6y�
 �!�+w�<p'���(�p @Ɓ�7^W7���	�S�H����s��x�Mv����}�� J���fSD�.�}�T�ҋ���7Z��O{dt�eg��:�(�s�s��˄���/�d�/N�j�:���Brb'��;]��}(��N���%�J�d���[lhy�".����*�4��&��&�����6OTJ��(����K�'h�X���UΌ�%R��I���]r�]#ߘt���v��|^�8�~���`�����s���a��\Ynb�J�9��g�'���٤8�����"��I[�^֯Ŋ�[%��D�d�~�*����5��.,�hh�>�-j����k^a ��7`���Iҫ�Pr;^ϰ���C�w�}�\r��0�O<xD#h�C\�<pd0������\���ɰ���}B����m���-��6��S�K;�ďPX�l��m��[$7Z>��԰�$0hw�;g^��/z��9�B,��8���.-Z\���!MH��y����	l
��9���p��>�q>����T��Ե¿i��ڇ�pD�	�Q
1�.APW��<�^t��t��V��e��Cb����������Q��LG�\��W:v�l8��[b8�l�@@ ��'��~���hUM�	�3a�-�ǻ���I�l���l�x�G�%��A�mq|�ުܘXު�\f����=�Ԥ��z腣ߪZE9�䛱!v���s��� ��^�aB��F9	h6���rLùyY��
J�Z�~娸k�BZ9���0�I8t:F����%H/Ĕ�ˇt����7'��$f�:u#�V{UP-�2;�r�l*r|h�(mV+� >�u��ˎA�����g�������[q:Nѓrp�&�Y���pcq^�Nx�[JR����4�D0�XqxCz#GY���Y�C?��p���x
�^Cs�Ƶ�\���u�|��A��]>o)
5V�r��S�i�l�\�a���
�\�b�B#�WdyM�W��P���cѻU������屻�v9f@�����C��{����u��-�#����w5�Et�Zo�XC���ط�4Ồ�|�{a�8I�!�Y䕞��C����Ѽ$�nyp��.I+d�*�$�N3ߩ�F���t���7i˘�삛b��{��`�!@��W�q�Uu�������,A�cP	��l�VFV�Pͱ��1u�;Cg�ED�,���x��8�m[4��{��w܃����n���]��hܽ��yd߳�y�j��F�EN�^R��0K��;�Q\��G����r�����	�8@�Aʺ����(�o[ŭ�z)��fͪ��0Ί���B��gNn>���ꕘ�,��w�i�0�(5W\zP�![5���١l��op�K���%��LH2�~�M���x���',ll����/
ڱ�`�×��s-�#�Z�:72%��S�3^�����m	
�m�4\�{����iM����6y-�+���RSu����tJ���:s�~"cݗ���ɼ%!9� �����;(�|��5<$U�
�Vv���5��Ř��=޷�E�ꖶ�Y�pB�b��py�{�5����\��Ծm�=����XL|BL�y�EM���mgJM.�o�"���x+���Qѭ(�E����W<{�}{#���O[A��|�P�-c��3�<Uc����.9�^I���(��E��Č�Xk"?��v'�-�z��9;�X1��j� ~��~k�lv���d�x�V̱L2 Ŋ\��8���S�1��IV*޴���yg�;��(
�2�c�e�����|K��S[��ێu��P��B�^>�
۵���v��&d����c�ަGϖ!�u(�[�����-fД���ɘ��v�аp�EM��H (����}R�ҟT�YB�.�|��` ��(���bY���M��IPI 	��<(ߑÿ���"r����̋�?�4n��t5�Ӫ�B��,C�~������;�h�r��.j���[t������k�'�p�vc�"�!�b�a���]p<(�ƍ�2��UeǸ�'�}�>G4حo���yCwv��ߗ6�n9��ȇ`2���<��j:/�v�p���n?^�:����3����՞`iH2ˍ�F�±�+�qI2ӡ��`�������p���kQ�����s�7Ӱ1�`k[b��4,/<v�a?�?@D�@4~J��z}�z�+AUX6Ҋ����/�F[{���EH-6䘯��'��m�TT�r�S���.��F�@ȃ��q*@�B�/�"�f�	��Ɔ�#6�R�N�a�h��4f1��7���dAخ*?Z��1�i#n��R.o<oA����jw�b�����cf�O��{��bϟ&SS���:��[̓7R���=�~ǘm�ɃU\w�q���Z�I���V�sȣG�#G���m�����㧔��?n�Z��~#�p��@�_��a~at9��\�C�_�z��ƃy�Q��e�E�/��p����������b;�h�H=���6�ph���sh��6�洪�ױ=�M�)]b�m�G�Ύ�������C�4G/	�C�����x�4qR,z�,�]�h�@ɠ�L?`�U�mзv*��%��{���N˙��$�w�H��{.{d%���1d��aeЦ^�2ծ��=���|s�󇒨�?��۴�i���<�>�15-��'$h��Fv�FK&�'�7�O��d��\z%bNיVװ�ՀcPԚ�{�أ�/
�֖/9ں��,
�_��[��n�(+/��OL�d([J�$R~R�=�9���$|�!�34�lJ�P/�z˝�I����/��'�-�e�~����&��ZD�&-����a��3AAT��䑛�4��сE��#݋Y�|��H���4��5N&������kW�Ԁ���2k�|��n��7(�q~�{�&��C�G����
^	?�:7w����?8I+7ǋQ�o��"�/:��2��>��H���2�Vf����<�!U������������Ci��Z*���,�(jc�և%B��Ȯ���>(��rġX�+'��`�x�������C�z���u]/�Ϗ��R1Q�?z�G(����Ҭ��CL��Ҡ�J����;�n�=F�˫���`gк�?P�ؑ���!�[Ga�T��3!��Cm���2V�Px��k�2���hP\+z?�������*�l�����D ]FG�)l!���a&ƶ�*�XWO 4Z"��*!�+CO���TDK$ɛ� �(t�#�Ai�Ɏ@�������|i{��K�3|$@��a_};}`���1 �ݖ���k�k}�Ԁ	��?)���5�xX�l
�l��6|��r�4~i�w�R�Q�·�z������\���X�@0��η|��:X���K�,�)�����?"55��=Pr�(Q Ʌ�_3�txQ�mK�+4�N�
v��� A��eF�.w~&��h씚������i_ܠ�T�ICӥ�����Vl���
G���X��ʣ^����Ј�u)���`�������ٖ���!�#o�&�y8���<�X�|�p������-*���Z?��6��~�:c�맽�^�EفiZꚉY�p����n��7<��k���H�ͳ�p���c��rN_n����(��#%,��"8VN�,nG&�� R��ؕ�Uc�1{;���澦�u2`hh�	�ڤ����v>hu�.����#��C����J
�m���/ނ�G��)P�Q�(@�˔N�����[3�+2	x+�>�ӆ��Ko�$~r�b*!��6�3���b�U�oM����������:�=6g�=���j{bʡ��@�ue|�m77��ǎp�e�r����F22�V�s������_��I���T�d��6y�\�)�[a���9ٸ[��6�Bc�=k�MהjM#[��s��gZpV1X�2(8�����K[�z�8!G��a6R*m/Ӵ���z��G�K����P^ ��%L�D8�̘ި\3�mTX9[����[ ��P���ݝ�&�����u]YǬ�濉�n7"�D�� Sf�t�^��`ԣ���-<v��iyJ2
����"�+ /�<ز�����H��O4+{=_j�S��e�#]XŘ�ak�|ڡhE]A�ۂ��Mw:+԰rܧ����A�	��yV��A��0U��h#2rPKx�y&i��}][W
24��m|Ⱦ.J�E$XKc���3$��}愵ڪ�����-�૸�v5=7�d�M��EjГg$Q_R��҉&�o��.��
�<l��}6	[y�r�I~q����z���B �KⴉSz1k�A�!e-�O�/��L픮v�=S��r>�����_C����u�!��΍��u��H���}v���vH�p�W�@爯���'�����<�Oܯ��\����nN��mr�AH�fa7�F�j�W�/D	<rŴ4��8ʇ�Uf�Ft99-��r5@/?f$Yd��~.O�	�i�=��C��`S��1	�$���W��>�\�[�&1������۲ ���w��F�b��0����qZ!�L�O�All� .h� jX��^G��YhK�vfN��6���[������f@����wR�S�]WK�r�����4ξ�~�b0Ct�P�m������E��f�[`��3҉�P6� �F�tNm��������������p��C~����K�è��l'}����(R��>��ɯ^ȗs�{��� Ӊ:��'MD�R����+1uK��V��l��_θ�䝘��vV�{���_�m�����VN~Ҳ������}�y<���7��6��k9�P�}蕅�"l�L[^�
9���-��m�p��b�M���}.I5ϲ_��G��e����Y�G���e�4�Qn��K�tx���kcw����@ɔ1	E�@��y� ������.��FBD������
+��[#J�C��V���৆rk�r��D�Q�(�4VѶ[|U?x�c���'��=@8 �|1���$t���t�&�r�޵���� ���ۗ|k�p�?$�֬6N�n>�,HY���n��K�8�`��h�Wy���F�H�k�Z���s�������j6g,m46�+���h�Ĺ*�7>�r��cZ�PcQ�6���`��Y&{�d$6��ܹ�LR�<��g�'z�#z����X�.������V66�!3��[����s�ܡ�"�Iڊ�xrC����P!`��Х1���ͳ,7P���M��G�]��X�rK���㎡_xs��m��f�{�B���<���tQ���W�]��K-}��i�(˹����%�Z�Ƿ��e}�C�����Ԭ��&oIC[��t�%��0a���L�8㪨.�6�wxs�l )5:%wz�۲Cir��x�c�2�y����
���A�Ѳq��Ie~�4=:X3�l0L��B�]w~�ҏ����6�jH�K������iѮ�qa�j�)�ߑr͗d8���6�����X�A7_��#W��O��|k�c�ߺ�g��w#�&�*4 ;���	*�@6����+�� ��{S�}Ls�}�թ��g�Os��|bo��ո�V��?��X
2���֟Z�jn�թ�t+}-mS��	&	���E��#�6Oݾ�}�wN��<�� g��nն.}5WB�(���yEUt����+�m��B��4Ӣ�~���-��\8]HPh����9�{�H��V
H��ƨ�@�b�`Fh�j�3��I��5_��b�-f!<���U�=X��5���n_dĈu�%6�����|�\��v�2��x��f�Y$��Y);�-��e���^�{�H�g&�N�(=�{�L�:y�hyţ�s�sj���~UdTv�5�E������@eæ��ظ@��%���*jen�tr��q������wD���DI��['q��^����`��aӔ�L�F�����\�����;i���T��[�TS���)���#���\0EA>�nH����0gge��yy�c�w03p&/����@E,{<5~�l����9�݆���;��f+�����GH���<�v�\$j։x���qo�6Z�k!�>7\M�j��Z�>��ښ��"s��.����!�
�>����~��-� ����i
��k�CX���)�MŻs�W���w���KJ�%M���"nH�_>C&�����Gn�!~L�5���G>�s2V�^f���w��\���.
w=�5Bl���z�����6p�_���i:�{�z�OIo1syp�}ݱkF�6n�-��D�Q�p���1�H�յt&a ���?m��^Њv}k�r�P�l�����y����.Z̜*�����c(����4�,�Zbo��ȄK�z	u�B��>�_K5�N�9}���A�x����LE�F�)ڜ��4	l.x������14P2���^Pxf���Yw�bE�����"*�ON�"�c�����+�P�� ��	���g����e�:�8p�i��RAxiXM���2�$��q��3.QuT܏J���.�G�~��^�vU�1[���鲲-�C8��"�)v��A^���=�(�U�+o�Kn���2�����iW��n?�W�ͥ�L�>K��K.���:"|tQמ�mҒ�}%��i�#�CCڹ߶t��d���l�(5
�O�.r]t�E/�?^�Em���
7@���р�d�p��W(����MB6R��\Qik���y����䰢{�Q2S]RttRAI{��I�.�p�C�d������ฏMV�_n�9�~6�O_���ǛA5�#��$տMQ���ߎ�} �yo i��ֱ(f=64�f�H/ܣ���h�ݧ��%*� ,��.�I�l�hۗ%)�UL�Mﷄ�� H4'%�*�fd�F>��å#����,��YS��iz���1��=6�;�>V����������d`��Bh7�ȞZC;ro��=)0�kr�Jo�N� X��;qPJ0(��$�՟'��vu�8hߛz�p\�O��k,K�b�ghSYD�J�1k3�����շ[����±<�%�hG����t�zÊ�E\��op��Qŝ֗ݑQך�$ٞ��L�e�I�a[6��%
�`�n���k��[�N
�����E\ey�r���-'�S��S��ME�1Un��1 �)�v��p)�	��!����lo�R��\mĻInj�
�i���ՁMgx�j�gU�����ʆr�a4��I5*ן�z#*1�$uz#����:ßA<�� ����7�B�d��&J��/�� á�z�[t.���~'�{����*�Fps�o@s �
�Cr���5�oqo�!y���:s��;�J6�б��uQ%��i._�	��2��D�g��2'?@9�昸c�~�����d��"�F0�Ax�"G�M��j�
 ��,�?%a�]7�tk�_{�E��lR� �X��(U$ �s8�++�xP|$���E2B5������Ƌ����� �g�༬��n���G��7��}�(�YG����N�:ݭ��:�-����j�H�BQ��@I�t��^���0�p Gg�����}�oK���9C�[�-G!�0�2UQ��63e��\�`�v�r���=�5J����i�J���3/F��F�|�R����ۣ:�:n��L\U}�_w��;͜uHy.�#ԙ��"η6u���6Σ�>]�]��\�ʢA�� ��h[��7�`#Z
��[����T+P���,JrB7�x�'d{+X����K�O�/5��0��b�t�q��E/��2f_��EǄ@n*Ώ ���sC疟P5c�]�dSz(A�v<��DG�	�Zx3"]:S����+(9��Ex�ע�����A2�8��A�����/�w�`�W��YēG��}�ٖ��Ě]=�^=��ϞG�h?���&'�?�3�b�_v��5֙�kl�L*$���0��ޫ �6V\��y;�m�ZI	x��j�MKA?Ǳ�c�D%�Dړ��{hg����1�~�fd�����s]�@�ќtw�"rr|��Y�*�B1̠p��	Ǻ�n�/���˹\F�~��{TR��l�ʈ�HK cZ;�_)�U�����RpP�n����<�j.�YՊ��5A��Am��>m�L��x�í�����)_�C���2?_��RIԈ�Vc4��=d�/a���{���e��u{�I'��������{5�$|�J���ujM���'ē��*�(	���P��Q�ps���r'���vA��><	"�ƿڙ8�{>�y�k�o2��*����;����.����R�Q����C�>������l�e�l�~4�;,�K+D�3�Q�a�a���Y�Yv���]�(f��IC�9E�jI+����ʣ���kN�[��x���6
ڳ��B����@%�n��hEI�\��˷}��a?����t�$j����n����EC	�=e\m�؈c��9�3X���?0�,��x�����AH�˪��O*�_ٽG�A��z������4�P�:���#B�G�I�����R�F8��܌٦.Dn�'yj,�p�շYq�	Ӣb"N\�츮G�SwAw@n���LS[z��yy�[�Gν�.fė@���?�k��``�m}wR��wRt�V7ʵҺ^r�`�*� ��#7쒉zܔZ��S{4L�;宍=Sa�'U��

�&f!XJ>�g���eǄ	_����"�c]`4�K�h���%��h
£��o���	�>��2�dtpg�տ�Ã͔���u�� &�-⎶�ț2i��?��*�c�b� ϗ�{�|Rp��\-��m���9�,�a��"Û(h��/O�M�'�;Fdj#��j�V�1k+���7s�if_E�@}��2TT�
��P13��&�M\����,��� %��g�?r�~7'��S������wf/�����[�e�)�{�d�d �'�aQ
@lQ�$ ���7[ �0�.*[O�j)�ˊdlX	��|�����=���?��YXz �(ae����$�sG4ԗ�>l_s���X+tq1��p�ǚ3��=���b{�oR�i���oC�t��M�QPu�@���|���Z:U���~�@ؑB�`�`�g�E	�U�l��g|�4����)���.���(���qoA��Q~���:q�p� l�������K�4���T��c�֊t���E��ʺ=��~ܜI5H�����	�|�l��!���n�I��v#j�c"�0����C�uh̦����w��<� ��X~p���0��ݱ)�a��J��hDBG�8�e�2;i�>��a�vl?*:c��,��4a�G��rķ�;Yj�܍�c-��2=f|��Q�<����X�?�'u(�90�/�������kB�:L�p����M��w?7p��-���l�ZG�#z �F�X]􍫲ZU|S�o@k��F�/��iҺ�����yZ���d~��t�.Aqx4� 2Z�;�ؙ�N7�^_�_�x�9�7�(y�P� EO<RǸ>�2��WWk�Ӧ�9��߅i%(�fZN~}�'��P�i`��.Ǿx	/�����1R]Q��Q<V}�ic��<�@��]UiWW�Y��U��S��i?��I�i���{	�dT}P�msG!0�;4�K��5���:0�Ϗ�����������O,1� xf�����~'w��
O��t��g�*�S	0FWT������`�m���蓖�v���OƢ���<��9谂��ce�t���$J�>p�-o����֧�7	��h4�	��\��j��~���Y8�h����r�OL�1��'�]����8G�X:��u��~Yu=i5�
E�Ų|zd$8!6#v<8t�vc����mӕ��'�����=�~��LEZS3��J�A����-}fMH��ts�r�sx_�M��������f�%w|G�z���,�ɤ-K�]oJ�1���*�P}8��"�����D������$P���P�G;N����Rg`d8x��@�蹟��#���$����F/�V����R�{���L�|"�:q6Me��TT"ޟ��!c�v�������4>N1F��ť��֤&Js�R��R=�=@�T,�8I���4�HL0OV��Upy@g��X���)l5�q`���yy���r�(�d֏�akP��?�'C�S�͸��Ȱ֚������$\�ޓ�~{g{�р�1���
��+#��Ƿ×��LY �n�������v�K\'�������D��J{�Qo�,��8�.�I����S��=A�鏄�<���*ƪQ9�/�b��ϸ,�Z�˵ދP�K|��)_�������Gҷ�ym`�G����@	�KE;��lt���j�A{c%�gE��Q�v F�Yk�R=���������U��t���yE��G��뱏�2�\�K���齓[�$�-��,��j�/+��q>ҁ��ܿ%%��D���(�����ptwxH�w�F�-{07�z\؃�m�����R���!��k����(O�OP�@Tù�C�������=��1�����ˏ&Y�K�.��wh{���v�JHQpP�&⩆;[����%:b ���T�	�R]����S�cQ�5VKSܜfv���vE�h�zz����&J�0���^��Zq�r������/���'��ּB�Y�SQ���G��3��`Mɺ���悒n��<��v��z�q�YC�jw��
S���NV�r�ty2�'{*\�MUKK�ό���mi��PL�K�C�2�C��߿�8��>���`����!)��l��$K�&D(ǘ�/{�&O��㷺ǡ����p��	�3�+�误WsT�YE��������W����Ms~+`�u�K���=� ���O���0�^r둢�Ƒ�2��-���][���3d������6�O	BT��mT�]�w�������p���?q�#�HC�Pi����g��<���G�	л��|�ɷ�]>C�:Qf��;K!Ljۂ�!{�wN%��LD�W=���-�Zwg�1y9�4x�5oB#f���h7+	h���|sݺ���E�}���AZ�ՙM1B4X�H���������V��	�r��!6!;�¢�Q*��@��LL0Wv�^A��P/��2Z��n�hnF:RL��v�J�����6<x`�k���:)/#�v:F%�'J��Ja	�\���(L���"/>����_���l�*����i{�qx�DH�%;5�jq��$
.�Wa_X�t13O���}H?Q�	�{�.�Y w�O�Z��a`������Q�u�G��o�F�7R�}zȊ[�T0ϤM[�`/̦zem��ɔ�׷W��<heY,����@%y��d#��u�}���	FK�����D%���2=�S�� Ӹ���ܼ��6Y����''?{a�*�!�S�i������%|N@
~{԰�0E!6����q�ى�u��eP�7C��wv6��.�ķ�~��&o���ͽ�����>5�+�=|��a���v�r��{�HNNo�z뾚����rK�P���O2?�� �!`��7Ͻ����k�2�f˒��#=�o����Ϩ�Ϊ���喝���d+�:7�b%JL
�@߯ᷕg��b����<1��݀�b*�z}X}�?��7�	3!�{�F�\��zbھw���F�NS��$�8�UP%�Zޢ�=3�O��w�L/s�	6�J�u��棯7A���-S��'����)Qi��UĂS,Y�+���{������_q��Ԡ�ڣ���|�\jCHB`.��|��m�)N��K's��kX�\�&�x	z���x�&H��K�{=i^��ي/w�.�/)uW�-$�P�7��Gc2ښ�Կ;�Hv����iⴄ:��`�T�"fO���g{�)�c9��?�vg�<�"�j<���r&�����0bCE�BE�1����h��a����;�<s+BhlG�@kD٨l
���A~�����ۧ�r8���_k�4��3O$pp���1���I�8QqQ�XY�;��ń��A���z�WV����~��B~��#Ov���wC�?��U����@ b�y����m6M4�V|�t�����y���'h�tN���[l��������-�v��?�-�G:��[�JF�t�f�������开ְ�-�]�+ʥm��לu��ǯ�y���q�AV.��a��м7�˔?��<!@�����K�*�.�'�c�$�w�����8����5�2_���]�ݪP+�2|󼉛��'����;Ĭ;&�������o&�$�Ey��w>D���<j���(c��+�/	%1����[�# �������KQ��`���B<��8��DS2��Q�s�F�w���KJ:�����5.m:��@z@�#���p���zs]:o7�:�ϟ�b��ɇ9�:GI�`���{�\��dB䰈�Q���}�t��q�F=�ٹ]ļ��4`:��Ɉ���KN���F=>��V���vͷ�:i�#[H�=!V��b5���}҈EUK0��ٛ� ������U�r����֓X�����:9��'�e+���+e
��l��?՗*ER ���� kp����j?U�='�;shNB��IUee���1�
���oL��Ym�\���xxlĴW�ƤB�+��b���J�.�f蛵�%`cc[YW�yL�͞�vKȘ(L����!z�Ú3NC0iz������ETUk��7��b%@���d��p���dF����ttI�s���'��<��aČ���z�����;r[�	��b�G��T(}�p�n�ع���R%���!�q��@�Y����D����&
�s�:���,�{�ۙB��Ae��u�J��s�Ζ�ȷ��Kb�	��U.���./�������J��_zZ�Q�!�b��ڴe"ʽ�t��@���ż/ќ��s�~�?6_s���B�Sq��Db��=�7�+̰�-���|3WHvC$�<,����=ٔ�ퟪ
Tb����J��eD�1� c*������33ˤGX�FK���5��Td��Y�'͹����H��y~��C�����+Q��3�m<�:U��A�����C�+�5m��O���.4���UM�`���:�N\r���m��.�e�.���'�%I��q�i,����m!� �wM06�����J\֊鿄�±�J��Z��3�����9���	P'���:�
�Đ��*�<�dTht�R<[*�n�o�6�"�s�c�ވ=P��uG]�/�n�c�	����.1}t�{��"#�N�Ǿ]�&2֖@���֙�k����_Te�n	?fw���im��5PjX�C~Aeaf�.� m��k`���9�5P����L���-�����A���S7�T�A��2�o��c����"ҝ(�ok�/O������7���i��i�����^���͘Yy�\1�ϓ��~�4QR�1)-S+�nE�G�0�v�:i����$&Z~.�{�a�c��ļ�_��f+�c�?s��+��̊?҉F��z���UeiUY���w2]�	?r#|`��-��|fz�xsOئ[c	q�^6H�\m�����|�������l�Y�Ý�������C�Vu����5�k�/�J%����R��B�Vl�7@of*uq���a�C1�+p���=����C	���;c��Ŗ>�O���Rr�o�����3�4����eb�����I[�TZ������sE[�rN+QYuY��_^�3S?�q���*���=8�k�N�	��n�V>&��ѣ���� %E:
���-����*��"
YKR���Xe� lW�a���!�����t�� �c��)"�!��Nq~�;jE4�As�j�w��YՑ��*��1ߚ�p{�F|��P0L�jES�` �+r����|�������BP��� 2��Ѩ6���@��7?�o�������3�FyZvA1�������h5�����E�>��2���Me,�BHjZR��J`��1�WE�^� "����Y���8Ơ�{dT��x5��oiY�V�҆�}\5;��W���̍�g��6�0%��ja4��x��c��`���y1��2���Sh��V�����v���P=��'�^��w]��t:oi��4��=�g����E�#4�����u���%���v��Wo���l�b�h>3���AW��yHrj����쉪3�wwd�all`�
�0!T�����L�^�\�.�F����b(u������@�N�D�(!���F�o�q 粖��.�Sw0N��$��)G.�?�E�DX�Y�iV����Wc��n��H,��Q�>𩑎���*d���0jeO~������>���a�A���r�lt�N�#9��n�|��MѸt', �0�>��S����Q��v������	�"�.<�9��-N!���N�Y�>��V��y�r�}yEm�^뇣���j�H�Y��:%���`p^�0���}x�3��u��)!��߇;ͨ�(���~��|t��er�]��|06|F�/5�	y�:!Ho�&��ޥ�3�pL�����"�?���!�Y����[~+��E��p5��ݻ��$v�e��\F�S6��a��n	&��ejd��&KEj�Y�C$7T����[���d�/�
�~ˢ��
��e>�)�����~���K��Y�q"=�F�ƽ������0NⳣĹ�s��m%��(-eDΙo��OTS��!��Rr�	{%�&�Y[G���W�+�߰\�����Ϋp��>���o�(����h�w,�K䊊D�*w��/bL��
���<#?Μ\��GYސB�8K}4*�Y�0�зAW��+^����+1'o����FiYГM�1!�͜�R��A�������Gr͍=Q��R��� ��M��H���wB���s\Q��c��9}D���v�^+�����}���D%�/���x@s�`�����e�lo@v{{�wq��}X� Կ���F�p�o_���w��(*��-�A+wk�k���爵�ĝ�S�7u�\
 �s#�?��;<�����	O��)�\ {����׆E=���OuQ�T6Kn��=�jn�a�<��]Ti.�nT翨lZWvw��q��P�fo��Uܨ��s�>�Sw�]g`��B��*U�H̹kt��"���m�o%s�2��t�@���s�O �!X�^�^0�i���mxtN���aYg�n� �k_j����U�=̭V��Y	<?a�ޔ����$fn�ʹ��\>?,`��o���{��>�dr���d�=��oc!][�:ZZk[��jSe,z�/Aۛ�k�� ��4�6��ϖ�������Z��~=
�ǌ�O�	?ӲV��.ƣ�����NM�ő\%9���
�_��L?�<��V�mdW�~W���3��i���p���Q_.҅�6m��l�_.�qlY��u�lX�f=\;��`�c�:	]�cbIF,�p���W�
�nV~x@�la��S*
�G��]="9�[_T�Lo����U7օ�����Ҡ��OB�@��l���Qq��XL��
W�>3��k�yݛ���>�����t�c��a��:���l����-]r�}�|����H�c�:�\��Ђ
{���t�?kd�ɭ�=Y�~6�ųH~�14K�j�S��>Ԧ��4=��06�Q�~u��,,��ѥ<�]Fz�����1�2r������Ý}�6H���l�<��>:�uGR�����R2n�yɌ���E�����t�ȅUc������g��6�䬗�m���'���ֵmϱ��QԘWW/�sͺq8��ip����j���s��ET�i�ƾA��pG���\[����r/˕� <,p8i5LZ��[Z�k@Y
*�c?z#0�鳞��V4+�]=I3��!�&\�x��~\���ϥ���-BDX��y�=�2jF=3^ 
�~�?�r]��,A�L�K>�&9�)d�����y���o��ɥ�`{�CÕ�|D�^�X-�o����d�Ջ:���o'��?����X���R!������<�54��)�iP���1�Cv�+0�o�x��<�&���5�H±d��4QS�� ���Kt�'�#���,��.{.^�}2��8P2�[7�����q�W0+r��Dm���b���U �"�+�uo��%�B�[ǒ��ڛ�'e�9?����J��X a�y��z�u��!����;yy�ny�ך��`G��l���+o�5���Gh�!��?J |q� }.
�������	ʹ������r���M%3����u�\$�(�o�''��iz|�B����LL��|��ۑ1q4,�J�/�0���A�i�[�}�a}"�.�X�������ɒ���x�e���H��$qPPB�!HbތE�b��3Sv�7iquu���zt���$�. �L�ܾ��)=9�KK���Y�㦗lmu�� �V�����Q���R��Kɻ9�@����S��ٗۨd��[D�J�'n8w�~���������9����ݵ�,�Au��v�K�9��>2_�PzC�3��*Au��o�NM��z��<؂�髺�?�/�9.Q=O�<�`}���� �+�=.bR34��G�MnO�ӸxII����v�ͅ��Ö�Ӊ�ҙ�f�s**��
�\<�h�*2|'i�$1���)v?��$Ͷ'x�ğ��Z�����roZZx��ʏ�M<
�/(r���w{����9a�k���F;�'b����.�)���hi,�����G�����G=�;�.�/�
�DE5��>>b�3�kH~�E`z��E*E&�.G{Iס&�i.�>�o�V�88�dA0ti�l��/�c�y3�6([?�."����s�I��Ɨ`�}ϖ�]V�� ��Gg���u	9K�z��e$pP����K����X�Tޡ�fH�e��9��M��a.v�p�\��e�ӹ�GO��1�ZK��(*���U�P�����77������6���V��'��7����rG3$WE��O��Su�3m�f��������ꋇ1C��K��;R�UK�l�4��ԭx��l��4��Z:?�-A������O��O�%�s�K"�T��- �!�G�A��fL�3�����{�u��ۡM�~�zð1�Q:L<8�<dw�CPmQ������SQD�v�Fz�y
-�u��:�E���\=osh��n(�W)~�i��=��\ov;�~�a)�r�\�DaE��J�9�D<�����A$�(T�@�^�!e-���������6���O��NaX�iw/7EvJʵ���SGO���&����l/�����f���Z��T�+�߀�9�Wy�j�*�u��������Q�K�E�#_�]�����"�
���#%�{�b٥
o)W�^�fw�6,>b�qog�0���K���L��QC�},�gm�U�?�;�:)�LEŹ����a�����}W��Ŵ�N�R9��>3bIŅ����	a�/�s��vm7cA�K���ä�4x~�o�
�j����ъp�������6��rrn���{��f�l�z�S��$�L�G��A��Lqָߡ����eUTf�����6�f�i)ŋ�"mq�)P�whq hq/�N����xq	� E��"�|�y�{����ʕkgwfg~#����=���n�O�����=ǓdS�N�B�S�#[)�`�A�a�<my�g�!O%0VgI�N��O��#�/z����U/:rD�(�K�N���k�VQ����SwRO�����7��VI�������O�u���0���$
d�J�����Y��#�=��}��߆	�zІ�YA7ǀ"��[!����}��#ڮB�+h����e9Z����$���=;�D���>�vnX�Hb����J��д�x���c���D������2��O]��i6��.n4B}kb����;Ug����\9��V���Y��t�~�&p_`���P�c(4O<=a�A���[�潓P���ugyCMC�y�F��w��Q�����/�y�X�ñ�4.}�K�<�w����0�v�ܼ�W��?T��0O�7� R���h�-u���U^ЖBo���0t�lX<��B�,*�JR����~��&3j�nA����<���̥��������A!�t<�H0�.�E/�%)���S���<�~���;B���ƮV�9Q�x�p.�m�	��w���<�U<�*6�}wv9�۞�zo�#V8�_���Q"f=��93ݓ�@��Tݫ�^�8���mf��?���+�!�1(3KC�D�/u��Ff����Qa�r���5ݬ�fcV���F�i������M۔�=h�(��$�rV�M�s�)K9	G�?�'L��?}%�hK�y���jC���8ů1ΕNvEĨ��t��d��񗽟�C�?��Ws��x��!���;��q� �@��񶪢����5��S����bٯ%��L�m O�_k^�>�cV9��v2bN*���DG�A#:׀�����s�i�S�j�5�փԾ��ڷ�`?�)�!4�p�� �| ��;��"�5����v�K��t�>����]X6s��GEc��$�A쭢C��Ih��z�5/�v���&A���v�3��ׄ5��b����ҩu�TFt�����p�����O����)���!�����	c|H��u7�ʛ����zn��F|J�����f�,�Y�%����a��j�����2�������V}�^r���U��3�E�.���IC��LP� � Ra-��?�:	Z� @�]���,(P��xsH⨚�R���fKUn��J�Lp 
��}A�{V��C��{(kw�\�*%q�����l�~�XR=��l�f��\�d�!�߾���TO�J��ƥ���FOϺ#���i�w�����dB�hŰLwx�觔)�D���5��ܮwZAO\L̘�n�)0�c���Z!�z�\��'�)S�qL�Y�D����ƶ!�^݊Xf��`y�l�˄�Qη�oٹX�ډ����-��>W�9�w�ew�}!��΃顡�uGY����ܗ�G�X��t�"=�*u⯷���cю�8���4�LK�xU�K�������GP�2��vKS.�i`M-���$B��F�#��)�������Gl�Bu���řwa��w1ܙ�x�|�  W�*���꽸?'�j��ts�+�9qq'�%
�V�&=;�^�\f��`a�Hz��η�L_���w!��Ix��'Bz���U��<'U.�4�v�A^7S����Q����cO����y��&��[����dES���G��5_��~=�%��X��󟚯����Ǭ�1��{��}9�zy&j�А���xU?���	-DO�?��T��Tg�1����s��.t4 a�`�}z ʒ	�H�w���F-�z��[��!�^�6DQLi8��pe��K�M+��R}ܧ�)�c����v���#2�J�A��N�G��3�(1�=ߙ���*$�9!q���[m6:��2|L�8�ƼmP�����+��?�,B��|������8��p��v�5��=-����MϤ��Q�%`�(�e�w�ޞ[�?|%�\���@�7Y���ĝ��bJ�LY��Ǩp��t��@@���D�S�s�Py��^R%�+�� ���.�7���5��(%a�O�}�y�I�r����`Hf��j��&�e+Đ�E̳�6��^�8��)��>i�uQ�ڭ[�-���6��(���x:��c$�o[����+��	7KN�W#�~<�[�N6YwU� d���Y5���!8c�w������?�??��(�ɿyR�O+�d0��wE(+٘]$}�wR)([2r[��,��
�kT/$\���}����_���f�Ȯ�nU��9!{�WSפ�g�i�<?�z��յvH$z�zR���AZ\O������������p�/�lQ/ճq�rs�(a]���`�<ȹ �4����`*=ꬢ���H q*"4�(�@�̢�G�<�=K%��x7m�?J#�%+�y�>v��=�Ӗ��і�96K��D�������(O`浺-���~;��	Zhі�iy+8_!��\������֗< ��m/cem��?�7�h����L���X?�~-�Z�nK>�5�g��<����Y{�yV`�mwS���]�-��,f^u�G�\��d������s���}���/H�#�5H�������}���O$�HKv��-;>o�	��9���5�[H��e%��4P2�bQ�Ι�Iδ"�[�o_y�����=��W}�u (�c��i�qr�
���!��������~x6j��#2��}#��I�5����|NI�i:���t,b�U���C�2-�NME���6La�K��T�8����}�sN��81��=c��U�����Sb�p�c�3z�B����)��0��Y�dv�b ����~�z2AO�
؈d[9���#UB��ח:���r�����	9#��߶���x3;�[0�(������T�q�W6�ˡ�+���2�|�`��;Ә =��Zު?���-)qI��J�>��<�E5�pgt�+�eš��yL���#IN,P���!%N��4��pN��]���K�q��~���D�x��5r��T��|�Fݼ��ACh��;�/;Y����`YDBo��bo	b�B��bv��I�Y����9�s@W�ƞ��t�Z��b-��M�D���3},����&t���;/|�N�e��{{��������OO#i(��нU�ɻ?$~�]�*JrRԊw��ҝ��6����y��Sz*�jxTg-w_��
���haXtd�h.n��y$bv-��մ�6��;��A��ڡ���j��Z�� ͗��}��;GՃ�~o�$�Čc����ǎ�N-�N�X�>��;��w1�OD'�h>X�W��3��E?,�Q;S.z��J|�y�Ct ���rd��E[Q�=�F3s�����(����qgt����'J��H@t����dX��R��dRf�m{��{���·���l�Zf\E����)��X������r�h�z�����}�M��C�j�X�?0����Xn�/`a�a��p�2�Bp��<8�����H0^&{��5��֭�'>ǿ����͈()qu�!C��ܑ!Kw�����7'�|��"��.BI)���K��ں��b���N<�HMU��4V�$����ѡ�:
�ftd�mM�;8p-���s�2���i�|���9S�xrU[�R�y¢������l`QpTk��aA<�6���,�K�;�L�k#�J���ØK��P0��Tf��1�q���D�Ff,Ȯu"
�eG��H���߇�k�'��bf�2��3/�����N����~*��|��IM,����]�ؕ���ɉ��������J��
1��b[�=e:Ժ���w^���܁VA5'�ݿE�L��C[����u-���(��Z��`x���,ĭ7Us���D�L\|���`J�K]��O�� ezi�пKwar����ב7rB���Y̷�z�ܐ&�׎{s��A��.�3U�j�@.�E�I>�Պn��||�gGm�΋��+�#�Q�t�)p�Z;'�y��|Z�r��Y��
��'U��o�ݧ�]�1��J/?�y��s1�T�Ro^M�1N�;?��_�sw�D��vʑ�mn�O��}�jU���ݮ��J[[�j�ƁΞ���,ZWz�O�j`���S�t�=%��=���I�!���\�AT.զ��\����^T�'��Es��rr�}ݢK�e0r$w���~,�F	�zg�\~7[��_o:���\��&�ޗ%�=S�K�J�#��o%6N>��N
��a�h��
���o�b�b�_�K���jALN�$�j �0��i]���VQ9RA�S���M�Y������Ԏl$����݌��/�(P��L��rV�u����9w��ӳ�>�*���x|XK�ٰ��]���~ u�����b'	���ɉ�Ãd��D��7ϊJ{-|!9XL�j2� %�E��a%��O����g��̖���	�X�}��ͽRf��� ا��b�>�4�e��x���Q�q��dN�ZX�?V�<�oXy�k8�½����k�f�{a�#ݢ�M�M؂��$�ɑ��\��n�i�2��Q�~�iyv�iʹ�w�G�_�l3�g�&@�ڱ�1�s����z�	I�"���p������ja#"�����q��6N�k�o fA$��>Ivfw��}7��,�������]��/��KQr�u=�[���<O�o�V +��D@{\�0[X�*��Uky9I���Ɩ�ξU4��##�ٲ���aʵ)�G��^�<0����.���i�E6� L�w�C�VD:@��a*�C���=gN�%�hU;l�㢞{��OM�{�;r���^��S��O�G�� yWuߖ/Q���c�;�ѵ��֗���y�S{���n!���0J� ��P�Ε�Ir�闺|*�����r�$�t�v�֌�������k �)�V�E�h�c�xv�O�*���J.����e�8w
�<�@"�q�O�w�Y�����ng�ڟ
��T֟�U�:$df���>��ɖ{���tOt�Pg^�������a�NH��H�}sE��;�m��9�(�@��x�n�Z�;�T�)$i������E��Ә�~���`J�药֧Y���2A��#��甉���H�-T�t�Exi�~���ف�-ƶy���!���Ӊ����h��X��k]z���-������s�j�G�&�L�:��D�Y�Fu��@�1��	��L��Ԍ���DIIW���$��LY��uP�h�+�/�c�j��J��n�I��={�+>��(p���N��ބ�]���Ѵ�/@bC��̧L���?�"�)��bJӲ�Op���B)������<�;�/���ħ���|���5�v6��"P�~ag������ �(G�@ju��"�_����!}��FU�n�W�*�[p��6��� �T6Tha�nخZ�O^=��P)x$����� 	�����⍮�J�����+q�<�:�o�,�	�K�+�ק�8��ag�$�����0��ڍt̛�����I�ʌ�@��
]�D�3�Fv`�_���񍦔�os���	����3NK�]ei)���x>���+�ɗ~�.�v�s�-n�7�c�],H`��ܵ�^���܊^B�"_K�Q5b6hA�����_oϔ�?�{�tj��,��h��,y0{,�!�UuW� 
CI�����h�����N�tcs5zw��O����}%���n>K-q����+�3�KV�k)�s;��?�5��麳ToG�k�˟d>b^��s�\�>M�"-{38tŜq�즞zL��>R=�|��Oɳ���t.?��d"��c$Fw����)�ͭsӵy�Q/iD���Tz=C�y(�F��P
z�Ed�����{�����k�ޯ��fT[�+�V2����(�)w��{Tڬ�F ��՘5w��CR-Y���1KBb��s,G�,d�����1���bg��<���Qm}N灣u!��Rt�!�t�s?�X#I�Y4��7@mn�c$�|jx�!^���Ȯ�RՅ�҃&�xm���۸�f�.�.����8']tD��ww6��Z�.q�YԌk�^��}0X+�:z*ɥ��m��.Wi\u�5I���r+>|����K��H03���[��`��(Ƒ�H�J9��m�mv	������	���p�b��q�ݓ��Yr1�Qۓa�0���wu������l��R��A=�Ӛkt���y{}6h��� u��O��c0�AUC	_�Ψ��=�w_$�禨`xB�T��#��(+����"�@��D�b\:��E�K�;g��q_��9Y6�y�����S��[�e�	%J��qUg:���+QJ��S@	q�N�^�D�2y�ڰ6��4?�Y/�V�s��^�$��E��Kc�� ��+�_��$w��_B��GὊ�'��av3�PږG�AB�z�5�S	h�7,��o�:h\��Z��	��ȡ�,	������lJ��3�*h"3�O$��XN�E��;��:Ū����JN����r7v���܏ӈȺlHXA�YI�g8H�s��tld騄>��ۅ�K&�jcs����a
WB_������c�1<_~��+�B���OwR� ���7�����{3ܥ����Jm>!�����&w]��L���=����c"��� ����w�٠Z�ў�OE�v��蹋v��xW�y�[�q��ֵ(����V���(��n2�,�y���)��/����T�>���sn�\&,�߃�]ݔ�Q9o^'�h�#M��y۩y�����-,����JL�ɹ\�:/Me�{�b,�?���8�[�/ѱ]���Nx�NA1p�ys8���ט}>��&��M]D��L�3���v�^�0CbF��뵑*+�,ɫY}�x���r
���um9�0��Q��<����O#��&����@�K�Ek�'��B�M�<���f�����0³�Hb�ߩJ;��]�Y,ܐ��6��?C(JF6'�=@بP��w��+����Tw�'��7��~�tls����WX)ݏb����fݜ����#N��;@�5V^9��~�x�&���)�\2�m�' �����?�+=�<��`Q\yD�N�`���K��(x3��g��n����wx^Ͽ��T|���D���w���H>F��!.��Q[�$jH!E�]G_o ��v�p��%R�����ܻw$�3Z7>{Qb�Me��%NO_D���F�+o��,z��ݰ��AQ�o87�F'��P�-Y���;'��(����8��֒�8̶�6��F��ZG�͖�y@��74�7c6��X�� 46Te-�w��������؜=T�0��w,7Zݿ�D͠h\���`�5ҹ=�'����B��OO���5jM�T����t�p2�;���OP���^A����|V�{�#��n=�-�d��$u*���3m��r�����<�1����9gI���;�A���^H+��w�j�2JU���CKns9��K�mWv�v�m
(?�z\5���_�E:E,�ʹ�;�(a� AW	����,X��;5Ĳ`�E��EG���촊-O��(�H�⋶	PFV��w��7��FG}W	I���(�Ts�:2.[t��~`����'}�a��&�ngbf����Þ����q���.�a����{R�#�������2=,v�8��%�nM�
�R�ٱ[H`&��7�����C��c�L+w?��ž��<�:
�ֵ�"U'�f���%���a��[�/�$g��~800�ز��ꭧ\t%���&�!�8� �R	>aˋ�W Y�-Us���b����7�sfiZX%bed�sobo�����R����>���1�\FJ�����8�ٯ���9�?���D](�,NV�o\��р���n��+A�)���K�=�k "J/�l�@�ЉgM�2�b�<���T�2���R��7�����q���k�Q�	��_L+'���|t:�VK}��U |��g��/�#�ď[W9�.c�ana���	�O/s���q��Y{��;��M�֓u=�š�9~�@I�@;-o��y�����oP���0�6zK���+����T�7��l���TU	���1sa�^����e�!��[���?M���U���쥒�"�_E�ts�d�y�	y-��71�7����+����MT� ���zW�����#��8���|��Փ��b��YBJ*���q�fR���V��rd�H�4�z��E�N��N�_�����yip#!~9^{*9��b� ��[�P���zN����g�8�c�-&	��&(8��x��o�R�����E��~H��q��-^3"f�
�貉 ��j��n#/gL������9�uF�ذ춷_vb��x�o��o��]�`��_3����l�������!��띙/��dW�W �#�꼤[!=�j��F���DkkW>DtD�W�kCj� �X��aX2+%(e<,�JO���RJ���ﻡja�d��>��<"Ҏ&c��_�ۇު���M|C5��vC�h�,�n�L�l&�q�i��jp�����s�Z�fٶJԱC��Epu���A�'�k�:��&�_A1�F��/.���;[����*�=Y4��*�N<���+�>�9\-5��C,~�rmyu�]�F)�n�&�P9l������c����.��QazÖg���与���B����3�=��B3�c�'�-n�鏏�2Pw���p|0���8���N��"�n]1����a�����<�w���K|e���RY!``��Q��ې���љ��������'N&h�A�fJ���W�K�Q��Su�uu�)Ӌ0�Ե���Y�,G2z�������M���e��q;�M��� L��<��r5��	53zF���>��X0���Ԟ��j8�6�@�-�]d܈���0��ȑa;�7���&���8&Α�vVVie�N�������v�@��{����;���ۛ	��p���^�c	�z������SNO������tl'H���R�r/����=}W>(֮-F�=vj�HR3�N����1���)�nO�8)�qg��&O��Y��� ynY�*6���°�E�3�'�� C�u���-��$,��~�wU����{��
;x��d[%>�X
�u-��%��a�y�*����w9��s=��|�ҍ26z��R7K]��L�{��i��Iأ��c�� ����cV�S��f��k�p?����(e�;bq4l}[M�T	u������ʶ)��h�
d��N�E��d	nl?�j_=�1��;�?��$%��"PTd�eF���tg*I�z��nW�i����X��2�[E58ȷ�{ަ}X���j$�������#J����&]�8�Ύ��sERDcVl�M\{���Z�����П�D��W�������D�~�Á�/_ �Σ�b�ǫ�ޓ�	4Z�w�<i�Z�<�u���i<��b�W�8�1nN
1���*��M��L�F#���vY]"L-�#�����PsY��|ԭ�ZV���E�Qh_�:8.<\AXN^n��
3VN�E�3ɲd�|�B��`���sCMKЛ"��BM�6<�0�[������X8dL{�u)�&v�P.*�ב�ru�p�ƫ5�g������#(�!�s�>�дR���
��2�C�����!i«i��9��!]�Q�#HXw�ׇ�j��Hk��w��e��\E���KN"�����E�rS����ю��gj�j�quuv���IG�g�J����H,��b�1=�*^�OC���jc��$\L�c�*����，�NXꉺ�{[���?杞U�᩵��+���;�ь$�5c�85eJ��7=�D�f��vm3��k~������_�S~1A���t�y������c���F��8��]p��Q���$J�n.�>s��n�6�Vq
󈎖�����x<DX����Q�F�/�,�t9(3w\ �]:>�u[�|Q�a���I��Tˀ�t�	.��}.1"����Z�D��L��3���9�=������(P��&cf��	�����EX>_N�]��c��h����C��x`��Qc�>�P�>:0֞�Gj�?�!Ǡۗ�l
�zl�P���t �|��HO��ZM������俑�l��	V�"��U:�&kI��Q�^��d(��7')r1�R{e�����6ybd$
�p9�I�蔓��856 �Ƚ|a��ʍ��ZY������0U�Bv��]�g��/N������!_��]�]A���V)�����:3n}���t�(V�!�
��\��Q|�V�i�.ԍ_"Ȉ�s�<6��0,��ai�n4�%N��Lϰ�ps�~w_�!ec��|���h�	��,ȡ� M.D]�(�Ds�rd_�5/�/~-�A�y�
_a3�f���X��qN�S���!����=�7�Ȍ�,e����q��>_ەW�إ�B�)�~�����/4t�z�JV�]�1}�s(I$TQ���1\��l1T��\�az�y�?kXQb�X� �+����;�p��m/߻�~���m��G �WZR�W}�4�Ѯ[V\��=���4b��3�\�����RO�)).ND1�=J ph-�;��M?w�s@�V�-��C�9X�SE �/V\n��]ܢ��6'�Ygg�c�9����Y;�v�������M}y�ӏ=>��"�_J�:K��lj�	q�z���gq��G�#�v�pO��12L�ޠ�"�\Տ�L��L��)(��{K�C܏2�	�5�[���7w&�Y���[f���,���l�p�Q+�N���lH�^�!�x$�s�=�YV{v.��!���.ֽ(����9S��ʘhZ��:Z[�U�z	�}$s�g��(���s��i��o��Rϭ�ɚ�����
�������6Y�SD������5�[�L֚��Nh����վϮ}9`�"�]8�+4�F�Ak�|Z�=����:�W�q^:�B���7�D�����7��O9����k{p������#���髶��u��#��nf}̀�鶟��9�a���$��JDW�6po���IW�7���c����1!�)�`��f�|���ؗ�@��t��]�6��h2��B�(����;�B'��	�->tJ��E��}*�ǩ:Y�Ә���b�D5
�}���8Y�g�#�B(��,�ĺ�E��!������AU�T���ٌN��G������$������j��L���{��k�<<��������e_�,�SRm���Ɔ+<��a���_��;����tѐȂc>q��T��!����n*y�J�+u�8՟�)����j\� C��Ў�-C|���KOZ��\�~��t�j����`�����ͰQ��������l�K��{3��KW���ڠ�r��	�֖�>�������jb���ƪSWG:B|i��|���+�e�ӇD?�[����ev�Ƅ|q�!Ci>�g@#��<\+RVVtݣ�*}{��N�"(}�2|]���	�## �oGk�Doo�#���,y���b��t������a+t��r�K�u�!�=��35���=���B��M5��*�?�^ߤj�����"�
��;}�k������#�/}�V0�M��BO'���N���� �zX�Z@u��03��ҳ^������得��ʦУ�	�5����^XY]�G��r�T�}�,ƪ���I.)Itlk'�>�7���Pv���j�o�^�	�7	��Ҡ�������$�?�E@�eyx��9���~]f�5k����kZa@Q�X9�����4�$\�}��$6F�3�9��)BU%!F���#��#�� �
YJ{�]_��������?񩾩MB���D�;�`�=�F�'BÕD��㪠�쥋�Ο�!�y��zi�uYg���$�am�j�%�=�#Kx[d�.�ԖV�jt�l�AR��H�\Ƅ64�pLo��� +���_����{hl��3f�N�T�!H���09�u"J���� ��o�:g�r�$��L؅q,�w������Q	�4���Ʃu�c�Ð!dz�̷|��S�5���k7�$b0�'.G����4l��������f��?�m��>���u��ֶKֿT�wʆ���о���]J�Gp��8����h�E��jf&�lx�EOQ�.�V��Ž�:��!�2��*0�!0]��oI<�{3���$$����]�컳=%A�M��+0��r�)��:ERfvQMd�J��ByRl67�0 8�����y��)\i|�;	]�qW+�W�sk,�{©y?-�5��N���dz��"oj}ӄ�ZK$�g�,z^��˩�iˎ�����{��/ۆ(D�[�d�b'�l�e0�,��������x.������<l ΐs���!NWw�<>u,�o�d?&@��.b���6��S�S�/�R@p�}vg�&YA���Mf3��M�/v@���K"j����bB���w{ݕ�����
�/ߎ/V@��ny0���>;Q��?�l�z�$�{w*�7�w��B��nq��W>5_����Ab�!�E/��_����"Kq��S��-e�n�~��H�:-f=kQ�^���a�_��N��>6>=Fm�l�U���?<�9��f/��֪�e'�M�O�z��(O`�tz��zpԗh���q���ׯ�g-a�<��N��d6�@���ܼ蕵�E2}��I�]�d���o�󎈶��\���=۽����.�6�5,�[�O8?Xzt��,��u^�k��u�<�+�����:��S��L�w�����!N|ǒ��TJ�.�6e�E�~�*��
ye>'�6:��{^l�h�L��t��L�]=@6�Q[v��Ȇ{��t	p�|ه��M(!��x���_���9�=��;`�������,[��e�E,�_,I>'&*(�������䯶�/Ԫ��yk>�l����暴��j}�)�\��j\q{���G�`��1�+lu��)ћFc~%��?GGGAEq��(e���Ѻ�I?�&��!���!1�}U�$K󃭋L������v�Sb���&q�eJ$���������d4&����>u���9�����('8_0A!6bH�)Ƈٟ��V��o�n>�Q�N.,����ݾ���l|�82���ˈ�����2�Rk��{�&V���Z�';�S��c�/8����ǐO�n�Uڌ���'[���ږ&�Wl�]��1Z%����W��4�X�H��Fd��ER��'C�Щʡv���#6��9�ӌz��Z��1qVɉ��%Y���}�n�v��q���a�gw��?%}=6�%���`���.�(<�N�V4�x�>�K�B��ܫ�-�D�L����v�W^��nG�-�'Kj�b���-ٖ ��#����C��ͼ�t�w5�1��;��e���qU�~���u=ݝ������^q2���u���"�TTr0��5����bT*d����&��2�w wt}w��+bp�m�Km����[��g*)Y瓶� tE�ڒ|�ft��]� ������y���҂�	��:3��O��Q�嫵s������K�	�Id�����c�6Yk�@
�E+�*\�7*8!� )dt�7�9��ӹ�N���GR�/�8u&b���*#�漌Jz���( �D��Sp��={�R�RPT�ɱ�!��b���<�݆�T�]z����`ؒ�}��h*�](�j$F���rC�Q�/��h�m�(�N|Vһ������u �:Aݬxo�U�GHݭ�RBb��a�f��V>ga�K�\��Q*V�(y��2��dN��Ҍ�Y����X�{���c�A��o�9`���Fie��N@QS���V�-�}��{6d�u<���K��S��l�������ΣA*�{`�/��'�5ɭz���gS4�3�F��r��f"����|0k������n�t�t���T�(<� ���dF��b��V�S>U&�����B!�u��Bf��С ��.��^���}�Q҃��⦔ڞ6�R����S�E��Ir4��Ǭy���ǡ�n|�w��aăS:�hhxehbWc��"��y���V�k#��}ªΉ����:�=X�'	�2�ϰ�А�'5p ��W [r��I'�	jmW=:���&z�6�=k�j!������H���o4x}r���B�&�l��`-�wz�&!#�Bovv�7����j��5'�$e��T�m7U1/��ph?@�e���i�y�����X�@ɯjB�쐮~]��I�f������������^u ��$�t)v�,v:�<��E�'J��%�6��ЏS�	��� hY�	��5ӱRu3�����:Ơ������h�|U86�dl�!�F���Ͼn�L��YsNq�f�*]c���J]����0�!��f���z���jp��č���|�&ҋ����Q�s�)U��x���]��|>�앭/I�UN�.Z��j�<8�xڪ�X�5_�"$&.j�t�����i��5����%![�c�CDTR�����i���j��G�;���P%�;���|)\AY��B}�����V�3��H]OK��������t��X��u�xNJ��!�8	y#���8��Ϊ���4��5�r�X](=��褢#�[���+�XA�4���Z���"nl@�1�w���������-�ho��|�Ny���!��n�&-QU��f{��G-����1��|Eŏ��Ц16����v��L�mb$~��_���^An5�|O#��7�^��8�5B�(�3 �������{��������"I�q(�TA
')��*@Tc�@#v����cÍl�i�x�s��H�B��&�vr'�R�"�笃��;���&贜@4>>ް��s'e\���I���T��=���I�e���
h�ku� �ɕxՄe��1'���L��k����ߵ�Ct�"����P�s�Fo&�a�1ځn�&Z��k.`�ve��U��Z��6���r�}3;����8�ĵ�lH���^DSK޴����M�>s#��4<ZX��7j\�q��n�n��S~&��+.���V�8�k/Fp�fq����b��:>���vI�H�� c���^�SX��p����E��]��E�m�|s.�o��}\v��&6��`��l,�)�	턫��O�X�>,,n�p��4r�����.��&v�|��M[U�x������@+��8z.�|V��̀{�.�RIM��_%DC�c'��Y
�n�߫���0Tt}3se�|�u/�Q���7��O��m~�����'���Z����	���v����ɵ�J�����4�RΦ,�P'P�{�T�,��:Kɪ Ř���b�����
h�:�MJ�2m|}{�!��ꨡp���-�)qߥ�)cj�[d���	�������~\��P����q�q�z�|��������C��Ql���1n7��z�];�`�>ǧN�X��d�븽Z瘔������ (v���[�\�H�$_N�������Ҽ�'P	�8��j��.���H|�n��L���r�a�V�n��
rv,[��)�'|�����u���v��8R_��<?8�t�y�� ��_^�R+FT�l�?R�B�r0�0(��u����f4���^��$(J�~`X�7<���\R��W�9��go�s�"PA3~���+��&�&�V,CUl�,{=�P�|�����G��a������z��w�7~�B���,-�N�-~������R�L;����
��6H�`��il_��O��LӸ�8��Ś��T�`)�O��Zj2�į��n�gJT^�bg/�?}�T�&c�˗�0n&���iyY�e	8a��|���(r���ئ6���i�hO����F��}��ע{^RBdOWa ������{� �]8|���%k�k���JD>t�]4��!Vfi�/�F]t�"h��@I��Z��jjzy�bޝ�b襫�[����3�����1! B���xvڨ��s��ryLR4�§�"� 3��VP��΀���}~��ʘ�������D�4����v���X������j� 7[h�x#��黖~O���l���RK���ŴcP-j��=e3�n����R��+ٹ�)(���,l0���AJ��'lcw�4 @��k˞�Y^n��R��M���Z0��d.���B���bW^�����%�����D�~����C��=\�}e�����p��� [S9ҷ�B��@���Dܷ^�&$p�4u��Q�ĵ�
�j��L��*����|�JY8K�u�e�c����&������(˾.w�:7"��^����#��~Nx*s$o�Y�+<���G�o��=��Mײ��� ~O�щI�}cE����+`oAf���3��U0񩅓vb2�ɨ�L��<�y��[G[m�E:�!Q�ݍN"��e��'A��B����]�����x2>\�:�(Z�5�*�s�U��0Mz�m��k��-���"6��%?a'Oo�eڑ���2�!-w²��B�#����s���_}t|�����Ő����ӎ���<Z������UM5̤���{���uo�!����d6U�S�����wQ��&Fb= ĳŏ����R5�x>�w䋮�؛���9��/���a^e�n~.�hq�iq�ҭF֝@0FP~���ͨ���M_W�tK����w����n�}�	��@\B���2����Nw.<����Z}zw��OU�	�<te�
&C���Z����n�wfw����Pd`��kn�!��`E�L;K��W|is��7�ٜ����;����T�0���j-~�&�7��2����c?�U�W�i����+�����V)xD6���ŉ1��b�祵�&˕w���s,N�;�U�5�h����p�O)�+��g��-����§7�K�(��f�X$�Y{b[ܸ|�r"[Nf�0���/J���>~۴�FS>n�0uH���x����y�b�X�7AE5\�c��w`�ܤ�>=|��N�m������oQ�����'L�v~u<��l���d[�KjjZ����S�-�ОӉ8|�Lw\Y��)�W\d*�.��}���21L	t���R��|T�*w;���c��4��$P�y��%k�9Zf��:�x�&�:��@���n.���Lw<���h���*���j�Ǆ�q�J�Z�����Y
kJ�_�h�6�YFQ��V��h�.צ�TIc8�7c�$���1����ֶJHt����xö�*+����~6��
�mA`�:���2��0����������U@��<	.�n{���}=6�\/��֦:Nʣ��)�j�+{�N>E�����%:4
+x���-��-�m����r�����ry��������lD�(DA��3��X��e%ַ[����0�}��EE�:j>F��p#�<��QG�S���
�e�l�����.��{�Za%n3!e��X!:�j�"�� y���hXoL쉼X�\�l���_~�oC5�n�1��)��
�\e�~Ǭ� �P@T�e"����O�	�C"\�L�$����-:�g<t�Ii�_�V�gm�����rl�������ֵ�Z���`�h۲�O�@~ ���߫c�-����TU��=ߑm\ߦ\܏�u�-	�6t�qҤMd��U��F��P4#���!!���4���MY̩BoC�q��x���Yk��G�+��e:jV����6>>��--��_t�;�,��BȞת��ݦ��%�]�\ P��/�饑 ꃸ"<�;��E��M�5��`��5P�rj'~�Z,�$�o��>,�C�]�������g� ?�vx���b�pvH����� ��c�;	%����}�e���[�R�l7��Vf��������.�qq�g74�^!��1߫�V��� ��oֽZ$���y�l�5 �(�\�E��1b~lD�%*e����DSέ����ԖG�&[!B6#p9%�6ƿ>����j&
�O���ʘ >���gx/�-��D��bQ66_�c����x�+��\p&�#��~7TdG��\��FV���l�L(��.��(���f[���ґ�,��a���f�����^���@��I�Oq��'�T��p%���P�t���&x�����!��'Ąc��2����ᗐP�����{\�V�ڴHC�W4�|�>%Q4"�U�R;����|B)j�� �����7V^?�;,�Y����J�x�F��f�������E�=�O$NuU�@�GNӇ���s����Z�U��K�O�G�r� C}<�A>8O������=�O�߉�Q��+ߺ�v{�"�����7٥2l��ģ ��.q�����o}\�o0{l��KJ��da�Ca�aR��o��ܩ/�D�of�L�@C�H�?WW痆�ܹ�>E�@o�·���U�����:���A���_'���7R|�Xd
�1�:���� ��t��m܃	|����;Ն�.�Y+ݸ��[c�42���>[x\{߳�24��{�@dA�$b�^9���!J�p-/��{hlݳs�/8�s�?3�.�(Q��N��5�Cs@v��T�-H�ۮ9��	��\��ǻ1��)���@���f��(DDl�-Bv�K{D�C��2n�=�uw_F>�:tr�d�/��.{��|�fH���Lp^�neK���_͌9w7��k.pvߎ����7�=q�o��l�	����y�C�֡j���fBN�9�<��v<�܇�o9�~�9-�����������6'>�Wejz��%�2��[��h�a�r�i���<���M>nK��j��ߨә�����)�옹��ܦt������p��{��m�X^�LX$�2}6G��S�S��^����	����F$$�KA%��	��<�$�N��0S��$�<�u�Ρ}��p���ŗ�8xO���)��A��b��s�|�0;���l��ͫ(�����=N���ޗ�O1quZ*��u��jEM�X򤋺\:\+tD��^�W�f�O�3��ܼ}�&�pQ�Ը����9?��%|���C�����ʝ�IŎ6;�9��a=q��-�ᡮ����:x=b�[�����������ہ�DC��k�  ~ ������+ُqo�4�V�M���=<��B��^u�t�KA�YH�{�y���N:�"�i�H^��s�y�9����y�$�%[���q�'czV=_��/���n�����cBP �A�<� cRI�A�����{�W
�Vny���R�6a��P�FE[�P麻�ﶆ�{�J#7�����Q:�Y>���lZ�h��y���57�V�P~-U����	�ȁ��Ln��L��OJ�7�b����b��<[x�4��#6k%إ4�Ȗ݌�ⲩ�K������g3q<�P��C���܉��I��̗���8eB���(���w��@2�@A?������j@'���£�N��pGͰ�ra�7�4�[��@pƺ�]���טڼ^��������HP��ϲ`�HHC^_��괨?{-Oծ�����k&�V��=>�e�`iT�d>��Bh!ڱ��U/z�a���:C|�A���p�-ڗ�;1����y �d���qf���h��ߨKj5���D���a���"4۠�V!U���xZ�>����6���ߏ���^	����AR��f!4��k����4Ct}���_��[Ԉc:n:'��D/�����*�w$��II�=��|���&/�#3� -�:���QU�\�M�����*'nK��v�mϲ`AK�T�=�^o�áKr��I�Cm.
����Éތ�r���[��/r�VS�$fn���]@О��@Ͳ�b��֘P)���i�O�A)k�Y�v��2ܬ��뇛{B
���C��(�<��:�t�0�5<�o���iZp�~k��g�_Jc�"�)3�^"B?�O]�md�@��>�h�y5��~��)q���݀e259l�L��3d��Z�]�c1���{{n+Z<��:�^Xi����[��L�h]����2b"�1�3���z���|C�x �ܳ�>$�Cd"����Iy؎
��W����,X[��7�iH��'�L��/5����	֕��%z4��0\<3���y�e�h�{`���#�r0}�6�tߜf���e����y2t�su�v!������N��bͩzFa��.g�	*��>:E o�!���|�W�o̓�)0�꫍U=^ �gˮ����wp܅�����?�3����n*���i{���M}Z���/�Dpb�Ӿ ކX�)of#�р��A�b���"��%���hC^�Z�yw��'+��Z*T�W��0?Է�k�/��h������}��P�s0m�S͠=߂���������w}�Qn��\T�٩��L��X��С1�-hW��;�2S��!�D9���  ���8�u v["�.:Y�K�7��eG��ݪ�ͷ��h���Ap�?l�?}gBag��F�|UǬ���Og	?_8�7����P�|g�M����yUIo���S~������Ar���s+�XdH�	D�W���[���;�3��I&��q�1a�<=��e��.mr�[��̣���h
v8]�B�x�$VRQg)��(�Y��Ɂ%[͌����X�Ǖ\��S�w`򻱆�/4�< _��x/�|��-K�&S��D�V��AV�O~�.������QK�8���Z�'5��[��*_���:��2���=���*J������J*��ϐC8!`�� �~��>�ÛEQ�1�'武����$fR	�l�2�pM�It1���7~��wݘ�3���B��^{>����e	jd90�Bt;���/�hO��$@.e�&��ӣ��g�s��ԯ)����������Z��'�DhWuC�����D���'�����RB٪��������!^�w֦<F�e�%�>�ݚEu,��$&"h�E�)���%��!*EΜQp�-��S�o���hp�f��=�����s'�?6��'|I�)���?ٚ���u�������m�GH�pV����z}�#!�vE�-N�堏�G0D�O������x\c�]�=��(�k��{P^�@����e\����en�e���{�@��\E���/�d���������4�!o�MˆW/���l8�DN�`��\�dp�[;�\�ӀL�*�����e�Ϝ��:X���#z7�u�����Ӛ�\�#��#[W�=���Np��Q�$�f'���n{,��!�E7J#����g�����c���=~�um�{Y?pF�zZ佞N���LѺ����V$�"��?rl�����r�ִ-��(�v �i����2�8RL(R��%ş�3��-p�u�ǰ�^(���8-���=kQ蹾A�i��Dl�i��ڤh��w���A�I������C�����F�����H��i./�uN��E�$\�+�/N`�2���wkN�
����)g��0�=�~[�k	��x�@��{�/zlW24�gWG�|�������,��&��l�w|���� j̵���x	_��{+���}�nIʎ9PS���6�ݶ��i�������;(�d���@����W��v�/�_M^�]y �����Io���z�O����Y]l�J�^9��h;#��b�T`o��ܿ���DV�q,���rvi�9��:'g�܄13�'�� GA�M���q~{��&�T���/�H��Ti(�#{�'N{��p�M4?� ��ԙł�|}����=���_�zhM�=q*H��r".��ɄPVQ���L��Ŭ+�j��i��-��$cE��O����&�T�i��Ae�Y>�����{�=���2�J;v͝T��CX߱�^��/����6w%�<Y�*O�S�
��1�_ZO�EXb7�,[ڼ'3-s�c�x�������抦�4��3Ҕ�3�����M�R�&�N|	�R��m}ك�IE��o�|��]tMIȔ��v��A�T�1j2��v��bs���D���9�QƛD!�*aO�T�h&�I�z/��F�̉J)(hm�q�'V�����{�Y�)xʯk|N��/>��gIw��J�n���WO΅��|�SsѰ�\�~!�$D�_��������r�=�=R�NY[��n�-�c��g�(��H��VmI�N{� ��[�ի��ě�I��<P�����k����q���
q�]ё�wp�Vڥ��L�t5飖�v�D�P)��E}(!���WKr����F;���
>�_Z�eR0�NH@_ӭ�Z���	���
NE����k�ؘ�!�p.����w��3U0F�����ƇF�40`�j�����L�"x�	�\2{�����$!]l����n{�*f������7�k��0�b3����:.���+�~L�[.0�_�+\��=dٝ�F�������n\6����N}��q�7�.��ZY�gYR�Q��|�i<s�y}���Ws�F�.��۳,�!��㢷C�R��6r�0�[�� �X��7�'���GI�L|��=ެ�D�b����}x�jbG��f��۾���-F�<�(ݱ�Wf����ޯ�o/�E�,/[q�K���� l�?�p`�O����$��qu�	%���O�a?9Qw�?x��+��j�ǵ��ۚ�`�朘@�/[�=�Lj:K�9s]!��E���Z"��:� K��"!DY'�&H��м�*�W��CG�`��>�F��t7ӻ�n����RoM�K�{�	��uC��s�|"�����@������444��f`--��Y'c2�N�5���@YF�4,Y� �es�oĿ�ۂ�L�Tɭ��9ԝKEH��߆��Kܖ��(0L�՟ئ뽌!"AG�=r�N�I@�,�����d9p������A���=Ԟ箢��u[ �!��M����Ӡ�Ҫ��Ge�'m�P�d�1	6�a�#܃������{���E��(�-�&�Q�����=��h+.��:��ԶpJI���>[��9\r$וk7d��7_|���b��ڋ�X�o��F'?D�iT"�rlb��ߵ}A1�����
����3{ 0g��1n�=԰_:g��6��se��FVv;�� �;�?�T��Y�����_X�C�k_�S���ǁ]QEч��Y)�����:�#	Đ��`1�����ɕ�$���tC�\>޺���h��W�g���E�Lt[���{<n���3v�+&�M�Xg6��W�敔� ���]X>M UA*�q�3���t�\EH4��J^��֩h�����9U�'uB��*� �-�O$�t|��Y%��\��#ɧ%�,�aD�J�J��_��oD��Uy|wT%�[b���`M���!yhP��HM�_���7E2���יH�;Rڔڿ`����J�nz{�J�;�b���Z�s7�w�[]���g���R(�0���G�����R��J�1+rvG�d��v-�O7খ�t3�*�f��z��Q�
7?�8G���J���Sj
~�OL��ҭ ���Ka�1� @���1��7����1y���������-#�rmt���������VE��5G5ܟƛ�cj
g8,y
�,��\�{ mt�6Nit��|�y�A$kC�.�NxY�n}rM������S׾�qa��a�,P?���V�Ι� *D����bRg"#`zf��CY��N��������}�Nl�Yh#g�������/�Z�~и�a8R�=���4����$��-�z������z��8�Lf�.�L4Խ���l�k�훐� 1�=~JE���T���K�b�ly�X�hT�>��',�����Xa��3ԅ��yN� e�M#�k���Sd(���y��2��;}���,~ǁ������!�Ý�R�Ӆ���|��[��	.]~p;Q��Ud4��o��c��=�캐lPm��Q����v���Z5�R�����?��bhŚ����-�ɵ	�����ɍ�HM��x;�U_Y���+���l�)_yLy������eQJ��+���q����l7����OM���q2��p���Ki�?�AC_��k����~�iO��
2}����<������}��3���u���G��DH��^��F�i'I����y��v���4M5�v	x���^%�J�M@��Q�&u�!dn�LP/&,\|Mz-L_(a+\5�R�3ɤ?���n��ot'���ڞ��5ݣ��MLwS���H�RX�f����=t�-��Uh*o�ٙ��V�������p�-�%��vP9�_r��n�a��>m����܂"u!��TFP��"�$#�h�Or�_:ې�/�$�-A��o�+@�u��+:qL���"�UF��:Z�3\@n�K�bp;V́�m�,},Gg�|��ǀf :|�e�%��A��t1Pmdi��b*�H�x}���k�fS�43G����!f�y=	{5��_����7cs�a�`��cqcD����7?��
��b���#� uw������[t��ʼ�*��I���1��M������4qE�	�����M �v�Ce���+ŧ�q�Z6z��cw��'3�n����S2a aB�e�<n"��e/̴>�J
D,�s�����O}�������MW�0t:�}�3/Y���e����YO	�2�K���-
Xo�Ro�5� ����Cp3~�����IQif[+
5�h$|h�G�1^�!�f�| ���?�)�r�����r� ����f�F��?El�"�^0���1�
�����h���~���P��BzF��a6���������uy=�[�u����3Mz�����m�Ǳ�Sf�oa o�6���w[]^���yY��^l�H]Р�Ö��/τ���>Z��Z���Tk[F�z���T�^CċΗ�ͳm��Q���2TQh�����]$���KWo�cU�B���<�%�IwG%���S��/AI�/���v����H�����_�����6�Q_[�r�����3�pb��8���4:�L�1�ȡ�#�� �r�l�1��,�V� �� /������_Ue�w�޹#�e��D��쪀�*��"$*��r
�8�E�~�ݜIwn!S�U���TCUoCN184"���i���˜�2MABz"�~�,xi����p7�%e�R���"��e��y0;��`�
8\��%�)�O�*�\�]���75A����?�\~2�3���I[�d�+s1�U���at��_ȩ4�����i�k�66������yL<�J�Dʬ�y�=� �{<p�%�)I���j(&��ږ������_N6�d����,\�c�e&���}3���9��۽�6qi�,��j��j�V�c1Z�9�+X��gr���n�$�\���5\vc��T����X�A��D�Bn���t#O~�Pͼ��ӧh��r2L�Qr[0�F*�h�ߕ��{��7Ǟ�k���6RQyq(fl.丧ꖋ3^Nπ����.,Ƚ1�RT-D�|H�%0�k�4mH��.��v�;&o��+.�׷*�(�qA�����XD�j�'7R��/����P6h��6�K���ax�y~ʓ�3��"t��D$�?�+����l��n�����)�oam�ٴ+l����H�~vW�$�m�c�m��J�aǢ"��=���mꎰ�Pp������޷��[����}�w�t�ţ��'FS��`]L�d�v��~ŵJ�I⛺_���4���������0a-y���T@��?ۈ�/���n�y�6��6�QSu�Z���(73����w�kp�& .�g�N8�fC��j�!��� Js���U��h�"J)�Z<Y�i!��R�%O���	L�J۝�{O�ڨ�Ve7��EX���s`3?g���K�
�7�ʆ�z���X�����X���#,�� ��3��L�&�!�cXt�SMNr�x�G���9:�	�Ƹ����"��4�� B��[�X�<cg����?�[��ˬ�%����O�hR��n��*��7�������e"�u��ލ)�"�8=S�+�8� ����#}]��)�OG�H[�*����SX���W�2��,�r��l�SEkBZ�,E|�b*E�p�/��)�DX�'�B('!�ek�.���7�!�����B�1��~�x�$�%�>Ώ�5��>K�VΦ"f�ZG{��VX��*�s��1%q~����A�nS�ENvr�8<���п?p�W�
4�%����!	�|3Ĝ8�i��6n3a���Z������=���'�q2tj�B�s�S�EM�A��uw�������*�>���m$`��B�1<�N�Ʉ�����8��0�/m���<d�"�zw�u�%�>���S�M��:���n ��#�2�|c�C���/��y��ƫI%��?� �����Ē��D`R0@ �BW �hb+���`Fx�Ѥ�)��W3�O�ڏ���2�g��
d�i�.7���-׶q����/}*�{b��I@�E�k���6ڙ�	�b0�Ư��6�4e;��e����ά��1u܂'�ql��脄�����=�&�F�;m$9�rj����Ǚz_b�k���������1~�u@FCo��[��^뢺���z�ɇ����ek�j��(~�/����l�7�l�b��z�����+���v�$|��!1���m(m�Qe+9�:~ʌ��M�'~��޸gz�:�m�m�Q>�����$)�YV�56p�A"~������J�,���r�OCx�?@TAm���P���äu�6�9�Jj�`��&pI�^--1;���{"�5���3�K�E���Z�l �/�g��J���Q����������6ˎ��I!�u媴�+�4��q��/�܈�C��|gK{&�77�����Zx��)�7eg���^��/{��X0�&���_SWY~m�2+�٩�������m��-B��[��qaz�tE\�ǐ!f���{ǦrMp`���'���H�%+�M��U�߽��y��p��OYIT8a7s�e����SCt��#��	cfy�?}z��蠈�'Ej�đ��wKb꤂���^�TX2)�H�yb��d��g��E���v���@j_p��Νh=�W�D��M��WGk�3��?��1B��U|6Gt���or������	���Ҭ�������c�X�~tj�{i>�i<a�!s�zJ�DM9d�R��Ubq��Q����Y��V�j�R�!�%�U����d�H���\���J���f{��*a�U(ʈx� i]�j�
��y��a'2����A�����e�`낭h�h��2���L]�6Ǯ�*	)�gl8��}l2�ƦfX˛-T��D��b��1QhF�h�����(�B�>����
t���O��l?d(����ѯ�D�݊�*+;M()�\�WU�5A�z�����T��t�o��յK�G�~W��`���J���Ȟ�{��������G��H��{hl��}f�	�~��;�S#� �E\�LA���x�6olbwj-�q)��C������,�L�Py����5�r>j�L\2ȗ̅��M�����f$a�ca��I�*���_�ՍS�����)�Q9ܯ�#c[_)Z�\��Oi�0�w��\ίc�l�O6.0�sf�c�W^���Ą���`�vr������j�!�S�hG)�󫢺�]<߁273s�K2��I"y]m��ms�P�*]�����	��b.N�My}a��[�L�zX����ng�RX��H��?ll�ͥ��<��f�Sr��T��UBvZCAa�뙰�&�v1�s]�8c�<��J\�7�8:�T���w�bxKwp-9��o=���uX"8ә��e
�S�
j�v���C���<�"lؘ`sNX�E��-��'{f��^�h�F���=�ՎG��=����YFG��[��f��844uU��Ǭ���zWA��9��
�;����Xֱ�o�Pev-�Y���@�K�t#G8m쟏�x{e�p�1܋����{��e9y��'�n7!L=a�	Phr!�Ҟu�.�~���|b��7^�^��\�.LNS��A���:󘟒e� ��IԦoP�(Q���^��~k��=}=���tCׇ�Wi�TI��C�L�[H��x*�r-�6#ҀG�3���LM3��r�P����w�%vN�z8��X�ޏ�g���g:�7�-`L��,�,D�V��i��k��>�Б|X`����>����k���I�_�3W��ȶ=����������M�sS��Aq�?'5&�!���Y�w�=�+�j0���y{-�`��vJ�b¤�1O�Ͼ)�;�y�d1f.j���N��ID5�I� j�ߨV�h%���+С���<�0Yoς�xG˵u#�z���^GԆ��j�"��k6��mn1��j�� ��O�SX#�hI��"](C�*��u����GM��s�'���#�����,��]*a���Yo�]Mxo �&ݻ9��i�%3������m)<$\g�Q�-~|�:�n�w(�5���W�#���)3�쌪�~x�*��5`;ge.���~�l�Xl��?Hgn>v���::,="��n:%�� �4 #G��i��$�0VW�L|�o�;�|�'��X� ޝ�}��D$jg��_���QI7E}E.#&��l��;��l��#��";�T�ϐ�����@7��}�s���<#����Z��r
!���W�؝��=.� �m�8s�I$�J�Zq7�0d�gA$�"Z�n�ɀ�mA6�"϶���i�k<��#�8_�P�n@�<XpCr�t�����#*I����Ox������u�	m����Z>k�~�{��'�'S
5M8�@�o$�n�H�C��He����`����˴1�d]彞�'<���X�
�*(�o\oư���%M�ڟ�����r|�|��-V� L{�_�0/�ս���#'�f
�8-��u�P�v��I�S�MQG�0w����2�	fc��nX��#UM�n-����f~S8�x�������u�=���ދx�����1��ݐ�2TL*�@�&��3e)נ���K}1�\�E}��ڹo��
K`5?���Cf�ᙔ�õ�C���ͯ�r�_s��^p���}`'�� 8����]�=6�~���;�=�$�(C��C���	)���j}ڶ�.O�0�O��⪪y�(+��D=]s�
��n���P��ݣ�m��梆�	}�rT�G���8a����R�@�3��~�0kj��6]����[�D�r�M6��>����(�tNY�n�bЬ�mi�
'�	�&��kϴ)+��j�p.y|��d����Y��`��#���a}���YX%g�ܱ�4r�މ�ZCI��:}�k����۶�;:���1��3H�8�� S�-�jn.�.ɟ� �@����?�a�0����:���!�jf�3�	�KK@�� �^Eg?]���0_ў	(�����1�O9���}M�˸���>�ќ���W.9sj6|�2Z_���d�o�� ��_O��~Z�^s��f�k)qBR�0F�����kX�a�H~���.��|�҄�l���d^lW���Z�ʿ�)���(U5���P/a�ſ�������zm�	��ٲ��5�,����� ���%�6�����*���m#����p䫪���=#xOj�5����,�8"�'+�gU�������0lA>��B��̜�L�F��;���\Vf����-S��R�D�aE�����L^cUO�25?2Pj���~vq��4FVzq44>����Ͳ[��?]u"�w���$��!~�'H��E@��^u�Y�o2����~6Eo���D$����}ݭ�\1C��Rm�C���w���!��?�
�[B�G-��� ��n�F��'z֑��*A���k$�͆���q@���g�DK>Xʋ'�-�ug�#l?WZy��	7X8�>���s��l��/�{q;e������p��/�=ןW
�-˶`�n�D������k�"�%�<��jR����;���vu�(�0�y-�m�a@ĥ��:l��J3v}C����%�	ÐSB��l$u�T�y�&=�-i����gԙ	fzz��?+-L�^3ըkk��[�UqE��x�������rY�q�T�6�43M�b9מ�c�B����YXԂ����3�#���c����O��T���z@h�J���:��V"U�n��8�a�<�`�r��{$�a��^�'f@�l)5;�jl��k�is��ڳ������Jo�N�Q�(v���=�,�B��׷���>~��? �~
:�>MQ��Urq�o�\1#()�F���Rć��S�*��y[R2���_W:��+k?����=\!�U�[�M�@����l��z���s��ܭC����%��d��V/�īp��P5��ҏ�g�	�kLzK�c^�Q�~��G��W�	(�:�_bC1��h�8g&��)o~t!IL�y:4���������c_�_���W,�G�9~Vr�4�c�j�8�E�����Vs$�X!�����C�X6/Ɋ�G����J�G�S!�bΔs��%|�^yix:*�q5�3	J�
,���Y��}������rn}O���{���6����=��]�O��pDȔZMvM��YI��9X�ލ�M�_��&PI�����ict�����y^���9&ǙjU$�����bA��%�B�����݈�R�d*�MrF�x�(�b��0һ��/��lu�"�^Hi����ж"^�9�^���\�Gh1�ԇ����%g�E"���%�7	=z�D;M��(�.��@ˏO����6ö�*	�:����i������E�ux���g�����]�87�>���1��[��HR�z�O�<�t7�����4��k��D�ī��G�B~�(�y\����)��ĒiC�"Rw��������^&J��i	�����x���;Qa|�[(2���^S�>�=�!�ކ��`��}/r��$F�'k�Ye~9�@�Ua�X��/M��82�f��p����޲X�o2���&]M\�+l�W?��'��LYG=�ߣ�߷<�+c�c��)��G;k����L)�X�z6�x��W��"��#���G���c���.U7_�gC�0�Q�"4+������a9R�y.&��:�%F-�� ��j�K>A�����:]6u����&!�h���>��_���$�����s� G��u��3X�Ɉ������n.�w:�u�Y��DXN�N7uVy�\�i��O��̿�+����)���&μ>�p�K��a9�U-���Nj6��&O/��"=��ݐj���uQ+��<��O�����9c�_M\^�E�T�@W=�0���㿃_<u��NC3h:����*������ۦ�.��a��O��
$K%�3�����k�%�~��}�ޚ�Za�`Td��^U.m��N���kV��(��ϱ�/�Xg���>���>�����( 8;}�2d(����"���j6���R'�].d�WرB?!�1�Xֆ��dr���^5mtE��D�@����>d:tK��K�٪�+^�D l�V��)O�IZЄ�&�&"U���}�ϗe���zC��DE��t�-]ޯ�-W��J��[�l.�����}��EN���q)#�n���S}����b��>�,�YJ������1*'s$��B�}�&�"�@c�<R��51~�¬�|��:�k��.�sl���n��vq����?iy�n���n�Jc�4���Mf��	{1�͘� P�?�΢�e����A�BK��-�9���T{� �;Ly���E����=�D~�����5�oV���gt��]��)D���$�Y���(y�uK���@ ����5���Qh*��	�l�>A�Fbr��́P�!���b�n�iP��C.8��}"��C�I����,�� �Մ}���U�
�ە��Z�,�	�s:(������r	�?{���׀�+Ъ}v����yծ��/s���g<�u�����?�&G��3��o)�.�!�{s9ER<��A/;�iD�+��ÅV�����������(��b���]�������6I���_���{|�[z*1y:/Y*b��Dv-��pj7���Ā�/��W�
����˨;��.!���~7N�]��,qH{!QPc��M?��el�w����Yz��yd˚�����n���٤�Ӣ��rj�0�K7d&����� {�3R6���[-���-t#/���%ѽ�� ��&�Q����+ƀ��,�m �Xy���	�}�@}�o]B�1�(݋��4N����F���[���Ġ#�<x�i�<{Ǵml��ywBax������.l��AN����@�-W倘cp�K��#Y�Ԏԏ|-���j}��P<Da���ۯdp3YK�S�Zlr��� V}��m�ȱ���t�+�{��>��o�����'�&�8�'�k[� �2a	3�E�e�Eξ��-㘋S���3%
�ݒ���0��-��zlR�n_�8A\��ڛ��O��MR�W,�rio�J �e��O,1�/fX9�<U_i$�`z;���O����~��^�&�!���W�4K�������6
�{�������*�_�!}H��C�b���V�z��ۼaS3]��2��%>O�"`s��lb��W�wԄۑ�j �l���2���}��&bߛ�>R��>^��?'�O���M�:�yi ��_����x�m��p�Ё���SQq3'��|�Rj�D�*�2�is�C�]O�ݼ�a̋�;ή��W�.�2��uŀ�$�ݢ���?�7�q�-u
�9�"u�a���sW3��Y_����L6��4@*������������?�3Ѯ�9��"��h)��o�����V��J	D"�_�F �aUGua�W�s���
.Ɖǡ�
O7��KCo� u8�f�α�$�i#Mo�B=:2*<�>S�Urץ7�X|˚˥�GC3AZ��m�,	ѭ0�@��'N�7��Ax<�ǣlj��h~WxU�)fb����tJ�����p,2���*��<�KYd3����m�3l�`=��
����� ����ޣl�D�!�3����@�]h����p�N���5�a\�s���)
R*fuῶ�Ռ�I��qM	k��#Ҫ��-���!�� �tww�]� �ҍt7]J#9��!1C��}�����=�=��>묽�9�5�Zx���n�;�0X}�c-�Dz��������Z���6≏�A@��os���5�����@o]�).��D:�uF�'T�/����>��C����f?:���Ș8𱾳H���,8k��uE�	��ۗ�����Et�Ů�b!��Z����5�i���`����� ]c�+�υ�CkH��zL������,�������JO�x)��x(�ATc�!�!��8G�jW,){�q�Sc&�ٷ"k��@���>AZдf���w�`L�cO̴������ο��&'���ۅ�h�B�-���j�~��>��!�J�	����P���x}�[��O.�rg"c�e�L���8��@G�Xf����h�J�[?�=-Z=�}�	Ѳ ԣg��.� #�	�c��T���6D�:Ut�}U:������P>�<m<��ǉ_7��)7��3L��=��'u.駫 �5��n�h#H��t��x5��S��ds�X���� 鮬�a�a�_��f��I?ȕ����I��-3������o��|_�q
���.�O�7�N�<?^T�m��i0sQ�B`>l��3�`���vH*�n�m_�����Y�Fe�\F�a����+��ʦ�G����S铜_�Aic�-+)��gp����A��@�^��4�����ǡjq�X�tu���PkR�����u���"w��������Y��u^zl��=/ *I��g�ZB���ג��pn?^���d7S��w?{����iq��KMV$�C�䉿�e���=�7k�Ʊ/�͍	R��܌�
�#�6#�"ŻE����):��֍��ǁq���Y�2V�Yw�d�~Q/{ץY�"�z�z�ޢ�޷)����/1+E<Љ���s�\�O��{��FBЌ��jc���Gr\�x�c[N�~�~#f����,떙�&л�#fI-S>��)�һ1v�-���	e�=��'��&`ܯ���O*�� fmE�Q;^M��$���a���;�������ь�N�U��h�������R�[��_67�"�k���G��������I�t�N&@�k��Z�o������.��7}��X-<- !���!sv;������2�/|u~"����<a,|GdI���B��f��/�p��؛>3��F�Ԍ�b����u20@��`�@�}Dz�J{�|P�������n.a��ɴK�gn���j�3���Gyc���,ơݴ�K�Z���}�N�|9�N����Q�����p��^�������ܬ���{�t���^�hK5�Ӭ���w%�W�eF�W*��w���D/㫥k�3/s�Y��O�ܷ��;w��ar�0��U��Ad�����}����%ك�ܮ������4+�w�i�D�x�w�N��׺F}�g/p����Ʒ�"7O谛���}��@,����iߛ���kB��i�J�u��ޠ��Q�y���!�8B��1��6yvF̥Bg�Ku��ȝq$E����ֶ�]��Pr��ӓ��L��QE��xD����@�ͽ8�y]XZ�JA�YG	���~=��0���5�����]�2���
?d�͑����s��)��5ZP��B���x����M���'�L� D>c�?����l�zF�q
19`���-���b��@�Q�ly~ �J��
Z"����<��K��zd����J�}]`��B�+}�otFHϿ�NX#� ޵����g㬋����0jjDʑ�t���O��cpG�,��r�W�y�~��3���"��А���c�П$����ĂP,U!�̢�g,��&��?r��j1g/Ι_|mt5�����,�����5��O����7X��&H�-��co�J%�H��a��E�xo�%�ߴ�L���E_���c�3eH�|��ă��=d���n�U����5�j����v�1aW����/���>`����)[~%�\y��K���굈��eC�y�I6r�DT�d�3�GM���2$�7�.?�2�x�������m�J%$%K�0�8�{f�'�_��*	���}̧pq���6�B~�eS\�А����T-��1�����C
����+0���DK��+�,�tբW@�7���o�SJ��]"�5V6�yv �ٕ�!y�sՅ��`K��I��Q�� �����l�3:{�/�P�P��[�]����4#�̀�������VJ(�����J���5��{׬[��y�����8��L�U�.��V���H��xf9��8K̜2�Ԟʪa�հ;��4��6/�������K��#B<����j\�e�����-	=#>J����Jgw��7π?�	+i�K�z~�M�(�K
�o��DY�t�V�'o��oj�b�ߊ]���_yL�R��� ���W�orx8��M����G�%��QYJ�`檅���
C�Z�Uxl�Y�XT��j��m=�%*ϝ�ܞU&w*�iY
�.uN�ʍ�\��qu��3������Ց�X3�ki)��ͪ��w�E�F�QW!��6�ܿ���fa~��d�b1�[���d|�m�D�!#?��~��'��/���lEN񐇹yL��&�'/����~�@�"(�������Q�R����5�n��v�׫�[�e&��r~��u�@�E�^W)��QR?�BJ�������'���Έ!񼍴��+N�\���K������ȵ��x)J��ׯ���#�{����^Ŵ��w޺x-�ڂ=��D�g�c�����w/�pxIA��O���p�#���x0t5�q����
�y�>�!�=��62��CO��cmb颕_r�N�r}��k �O��1:�ص�M�nr��ٗ�Iq��M�����%S\ic|bHT�s9���]q�K��q�`�������j.U_��:柶hvZw��j�a}����\��>��ǡ����	�c�V
��&�;f���K���'��Ը�JJ`�;oo��*�"˾ּllsn!s�Ə5J��q���,u�]ڋ��bm��qo=�o=�)=�~^7�����f��o����^�k"z~"����b�3&5����ƛ�vŝ.��89��Tƴ���������ɱ�Qnܵ��t�ΰl��H�f�"��d)ǃ9R)�[�h&���'�nV�ah�d<�-P����Vo�!��Ƣ�-�5/D�̻5��5��Y��fM�K/֗w���9N�Χis˼9��ʼ ��G���#��c��#�]S���P����N�40���v2~%��5|T��b.
���ǥ��c�!K�EW���*��� ��5��p��S�d���mS���G�T�h���1o��	����C[*����:�#�e��!�~U�g��]C��R}�o�rW��~��n�'��y�A�i�m;o�v8�6O�:\��߆���w�T��sR1�p��*�]���x�_M��ԇ��W'����4�Mđ��3�q~����M�x�1�k��mEn��؋�K_�/��<�X�!�7��_~(�Mbm�6XaD��%�s�u�򖐐�+t�r�e IT2O1ꇙ�4�������ZK#/0��uU'��(���_l�Ʉh�e���$��������=�~��\�.�N��2f��W�zM����04E�z�<�<h��!���	EtJ#x�P�`&���|�������\�$�c���^gJP���� k�y"!;���y�8-M�`���R��G��"!�4�B��m���sY�}������WU`@O8��;<ٖ�	$�e��0�ɨ ��|zCT��j��y
+���*˧�
N���7�� d�Ӽ�+����4*t{��1,	xD���gc����>?����kz:inGgrl��n%�d��`^�/U��q-v@,�������s1S�|{�Rox�t�Ϥ�?��f{?�����]VpZ��s'�xB�NW�t��d`���U&��1RG�+�I�2Ǣs���N)�G*�e"�y�����~����2���o�8�Q��f���J�.�WUR�zO����1�v��[�RȊ}�N����g�s��+7�T�z�/p6eP-v��]�����+��$3DB�H��ăE�F�b�|��51=�xV�f./��ֆ���5���(�d���Zs�i����N$v�E���]��8�"�й�����h)�H���k9Z���f��#�%'|P���>�W��ÅV"v��|M����ȷ+m�p�ŸYy!��c�N!r��4�$�ʺB��´ �!kED!']����@����\�H���	@d���gk�7��_-QK���_qӾ�2�1�,t8��s1MHl^��fC����ӻ��i~�O�r]a1��HsF3}�Z�ƒ�X�Dk���\�2h��r�̘�`áx�� �*W,&/Rw�����ؘXԗ�@Z��^k�W<l�Y����q%Kx�]|�E��Ќ�v�{�.�b�7��$mW"�����x0���;�rZx�h���}������s��q�oo#�s�܁E�8�!񸕕#򦄉K�m�g3����:���l�À���.�r6�ww�pB��FPA-���iЍ����|V�;�u�6u2�)~Q�g�ڻweCk�8w��b�lƓ1��F^��dc�9-&�n��b/X=����#�ŷOD�����5�3޿:қc-� ܢ,>�x!�z�=�jYZ�dֹ*��8�UkP9��i�^�_�VVF*C��6�O��U�L�>U�9�ҕN+Yc�:j�a�V���@D��jC�$��L]$1U�[���z&,��J�n��dϡ���k�$d@`���U��U	�e6
�"��!}p�����Դ˸ ��I��o<�"S�C������3Ka��x�� �����((d*��xY�E����^�o<3PW������t��|��j.���
��a*$��N����6:	�g�=Jd�\p m����s)��ɣ�d�O:��G�����!�-�DU7���E˹�5R��1Ȥ����U\h${������"gJk�*�kt"���x�A�Ɓ����0#��� ��O!U��.�����*�G#',��C�K�pfo���y!)�x����}}�N�e�m ������$R��X��Ǒ�ΐV���d�� ����t!�PU�pӟ�ݧz�6SOvZ�[cc�.v-A���K}�@�3+��wi����Ъ)��Y3�dC+��ў�9q��r�5��X��ӽ�u��u��@xBVKQ�+������y��w�ܗ��?m��/���?�E��~� :�N��^�FF��z�w�����t�&�ן���Ȅ����Ą��`a���-= ����p�6PP�X��X̻��s����d��X�o�Ի�$����F����d�O߽0�Q����)�Z���m�����~��S��M��'k����'����7��S6���k�a�����1Қ�~7�5^�}����e�����?kT�)��S�wZ`,�7�SVV�=Y�Z��X۪�Y�.�݌��['~2e8��h���d4!����,��@�It��ޫ�OŜy�l�A_�%~�;>u=12ἔR|����3 s�dg/�Y��S;XO��0�{P�B �o�V��:7Ӊ��t)���W�Fv��'��Z��ǀ��S�e�}xU�O���%��LB�a���|�(;�a+�z}#VB�X����vf+��ڰ���N�=7w�T�D����$I�M�*h\.q����B�f��ƞۂ�6n�i �23�ڔ��O��I�Z��xЃA��Y��p}QLFN����G�����(�穪�h�Ke(�eW׎��U^S~Í�Q���bh���l�o\�L��[J>~��A��	Et���Hp"I�s���
����ߧ*a���2NW�U��ѧw�ȷ&Up;+��h='�|��[=��i�2�&EF���u�I��r=�����(���_�r]\t�%�pW�چ�#������y�S�Rj��[oQ�|�*^쥜y&����T�I�q���9�1�${hV��Te�F<�SҨ*oS�����Y�6���7���Ter��� �O�5�I�	\e��n�O�#���Z�^�/Ǥ櫅Q��%�p�L�}����kY���Y~K'|L�L�]��⟘m�-zq���tI=���zV��ypC`��Y��&�w�⡾!����4pb����:sg�@3)�G�A~�!0�$b�=b�a[������P����yl���h�ݎ5Zv��|B�9��_F鍳N	O�t�jc|~���\#4h���h{�������P&9�>[Hwy���2DO�! �ѿ�s���`ӫ�ʬ%���F����r#}V�IE�;eZ��f�@��/#i�]���~&�W�� g�MK��EX�c����$��+V�WC?���̊Rx=���L��Fr���N!��߿�KZ�GQ(Jp?_��&b�,�`���&�Y�^�pPOu&E�<��~��c5[Q:�.�ʽ�~S%rTy����B��C�����`�-���oY�����{���ً�m-��n�C�O �W+=#�ِ����x����gR+�R�ƺyŧ����%��ƥ	N�}F:��sc�c��~p�
�	o>6w��Q-���\�z |@�i�pv��m��~WH����"�~7�z���
rU������Z�s@�*�z��`�1���62�=�^���zj��Y&^��(};F^s6����.ځ4���ʱ� �;��q�7^����?���LK���^����� TF��}�*vU���vW��Ւ���&J��.-4�z�9�Rm�L�����f��K\չy8�!��[��+9K�Dy�@�:N� �`��)m	���U����HO]����mG�W��kz���	�&Ud�d�+�qj��V\�N�-�1)��Kʱ��aC��}��q�&1k��9�f:D�NRR���"�4������E���&;=)	^�&e �0N�HiF�Ma=k��j:.��+�l7���w��䮚����>������L����ןu�bn�Q�yiF̦��V^>[�"�|%�5���c���F4�Gj����q����WD.!dL����6�yun�%{$O��:Wڵ�_�M$nRAX�d^	d��Y/k�Nf�w��م�	[\XjjvУg��*U�x2�n�;|.�A��͝j�j�\�C=�9&�1�6��'���ػ[�h���܄ ��ֳ��A��\�#+���z�Yy]Mǝ@�q�� �oy?<E����bE�g�v��~Ӝ4~YKOX.�������<jﶺ����wJ�/�#�����)�k���o�_�c9R<Kp��k1��C�
�fF�}e��J����M^E��+e+S~���ױ�*��L6=s���5���/�m��o:#3�x����*5���Y�C��^A����_}u�����B��*T~�2�0��ix\H-|ɝ�F�=�o>��{��`>��s3��d>�kxGW���l�>���b�<Q��x� ����ش2�ӔfcKиQ�E;��w���[��&��O���$at�O��:Bh���!�M37�3ο�i��4��a�����{�Mt��_ jFؗ ������O0[,�����b��S�޹��h?�;�9����!۝����	v��\H�2�Y���;�ʳ�r�Z�~�V'ú��,�H�{@�T��L��4h����$i����5A_�B�2��82i��G�@^������Ŋ���)��S���_��.�>�覨V��*l��U��*_�WBJ��f럫s��󥸪/z�㉤8��O0_�
U��Z��y�*.���i�{_��F���	\U��+��2�Pa��v��v���5Nˣ��)�[���{R�W�]��Wwjj�jP�ќ���V�!)sQlU��NS7M�e�њ~}�>c"���u��"�	/<?U�/1-˝6.�R��"��!�+��G]����ь��F��ٽ&��4~�'iɶ��9�T��%��iL���{���Er����Mdq�l��To?֍��Vֈ{i�0�p,���Bd;R	t�Qm�JR�*"X��˭�G�_�.0���Q<���tm�ެ��@�$e.>�v>�.����몃���lwZvLU
���	�����M�s�d�� �~��:�m����J��Ysx�[�v���c�[+��2c;'�p�§�G�>�-�#��Y\>u"�H=2�MS�8�t�
DA۹(y����.;,��Չ~W����C�c�昽�^{M�OT� ��Fj$u�A������H�6�!X��,���+��>����"!$�����!�AH"Da��":�;��*�s��Y�����~����Axi3WjX�M�83[m�ry��Qշ����=�eBW���;
N&A��r�Zy:���D?�+��-SB��=��7t��%U��~��T��SM����q����!��C[��Y�\0�l�Z�h�>rU�TH �Ґ�,�
����a@>.��MM�F��c���+b��8rt��[z�አ�_ּ�ȅ�TF���z�2l��u;h|�:�<��q��G1��_MW�4��?�!Ë��b��HЧ"`r �����I[c�+.ޫ����Y[W0��u�7!�tyhA)5
	R`���l�)�y?��c�>��/Q���CAb&���,�y�~�ӻHEF+*����ǸA���,��[W��Rѷ$I^��w��'V��1s@Q�$���_id�V���ٽG3=��!��x�w)�q!2F̚���85h����P}K"ǚF���V��|�#�Y�n�s A#_~�
01E��zk�����n=�_��e̬�������Y��g���~^�Q?��^d�[+%�\��}m�͑���p�i*	�wҌ��]
��E�u��������Y3qqq���~�3�4���6���R�M|�98������t��W����i�����u"�1�{~`MLt�rfJ��f_{��7ތ۽��&e��A�Ԛ���c) :*..�o'�u��E��N�/�9j�w�?���戠+���������ՆB��]T���s��IPXW��$n=x?o���{�a��lJv� ��a��x�?�E�_g�	��M=�-�f~�z%Λ���ǔ��`\!
�5����L�k�.���v�=�'���{��d�T��������ERm��V�:��-Bե�f���dy��_cK�~���gAa�f�/��-z�-Ί��k���if�.�b͟>����^UT�q�a���m��{�4���`S\��ծ�����{~��t��kN)h3�e\�9p����?;;;�=}�yw¥�A��Z����7� �R�s�����[��O�p��#�#�LqA�}|l�22.�m/���L���i/3U�V)��v�|>ꭚ�"��u�#������}:X��/��O��%!��v����©�Y�l��V�/'^P�2�3�����/��ʭ6�
�:g��:�`�߈�cA�V����-Ĳ���o�O��ɺ�'���[?�={��Տ�ӹ6���IF�J�T��oh~����D	�压�o����!���񟇭333E<;L�O��Wl{���9�I�j�������R����J��/�^����']��)��[#ү�Y����**+�˫w�0���/��kwذ�j�j@��/R�H�e5,�\�}f�"0	00n�Q`���>b�JS	=N~���~�m�>M4=���S�k}��`����@�D{�}���`So�[u�[ۺ��X���Z�*
%@]@G��q]���t�L����:t�2�`���M`���
Ǡ�89��^��������(*))+�����x˺H-�P�F���<t�XO����P6r"ھ�Z��h�s���[9C���i�ivm	Γ�#^`O�)=���<�����[׌EFƢ���\��#b"��௫>��������'���t!�j6�Oq���vUW�=����E�Տ����e��>5��WI�oqA,�Y���酿�OYZOGb�7����"�������fL���_C�RU0���ã�q����$�<1N�Q�8�|+��}�񛥖��wW\uU$�b(SǤ��~������a�qn��AU�M�����7VL��N"z܈�g�)�}�U<� vc�������ҥ�c�cxI�oW�÷#��<��H����l!���hF(�l�$�����C�2F�a�m^�|�i�$s�Q�{
��_��{�%����%���Y��8�9�����r0�
s,W[:�����y�#_G	m��ks�����@I� ء���:���? �7��ƀ��5��8�2��c�=�ϖ'[�1�I�E�V�>�(�Қ�P+ڈ@^��zc�@'�x{P���$�
���%��&}T��@���C�XBzܩ�BV� AU�k?r:}�@��o�
3u�EZ�c�G'ug*���]#��-�I�n�S���Qi���@�7#�o¯Ϛ�/���Х��CU�OB�,p~��%�Ғ�k���Y�6��:�{s�sG�����<_�}^tK� -k�|j_�,R�ƶ�� �|�g�`���s�,���K�C�uIj[o2�:�g���	_o<�}6���X��m ����p�~/�uv��L�Fˇ��������v'Q���J4��]ׂB�XN�#^h��P��Ǚ���m�_[���wDYDm.`K��JxFc2��o���S�V�~����f65p��{H��A�h��k~ֈ�j���dU�%B�����Y��W�����؛���R�����f�$ݏ�L�(�w�����͚�-�D4L�6w����ښ�I��߱xޓ���\
h��xu8�}oDg�FAF;)�Z3�v���g>e�9����3�~��TU��s\��N�e����R�^����Nt��t�
��]w������픎.�t��,F����Du�f��z�e��N�|��������՟g���2)�[W������7��[*�?0��!~�m���A�7p�1�G�����q�X���A$��^sֱպuժqf�t�a6h��I2D�khD,Βr�dC���vr{��
��<~.���Ⱥ��J�V6�;F
p��{��ZV��R�Q�|�<�w$�c:�r�������m>�%*r�����t��h�u�B�������nR?\	'����aG+�U[bKA?l=H��7ZM��ćCx�GE:��"�+mщ��������YuX?��R�;��k^;�أ?˷,RM����;�_o����^kx,)��UE)��*i��h�N���
�4�,��p��E���WN=����JX������e�����5@���iT��Q0s]r⺍�e;<�� ҂��gf�e���M�鹜�Gh�Y�e�8�Q0�,��":=�tvǇ����s1S��Y��{?:�����dA���lxS�99B�B��_�k˜w���)��/��N�G-�w�`P�l����à�I�q�+ʸq;�]��J)`�K�=B��h�����G<Ph/bK����]r##0�����^�����!J��gN�"���o��w�i��-�����`��ŸF��3"�:��
��/�S$�5�a;��͵14W�h���G��SB��6���%ƼI���7a�C�#�N觫T��A[�'rs����q�2R,C�F���B��(t�X.�^*ɣ�=�ޟ��'fQ۬��l��((?��;���[{8���9��%I]���������'��F=؛&���˧�-Ø�W�����rg�K�8�YVm��_C�q�j�����Xީ���#	Kc����-N�^%���y�F�v�nL�oM��&�ij!��3�m�r��8q��s�%����<�����.��t#���n6�\��z��>����с}ηU�G�2E��t�����]X�]z:�t�T��c�3�V�H�\L�i����
�����~bak��!�p��"��ǩ�^a8��eF�'`��z� ΃iݎ��1�̄l�	�U��I����O@�=�G��kǽ&.��͘���}c�vd�z���}�?E[5^[H؞��gcgy1�6��^��XS���U.�WU�(tFRO����3U��畷�����t�v|[��:(�@�=/oFo�#�lv�,�Z�"�s�[|m?�V/psR,���JF���÷x�woo�GJ��|�P��'38��	�!t'"�[eܣ?y�_��]��i���s`���o���PuA��}J�V�9�n�ܐ�Iw���x#E�`��EG1	���e<�k1�ᕺ����[��[�D��eL� ��3<�M���������﨤���:Y��}�� �vi���F4u[����r��bA`��:E�c�)%�BU����v��퍱m��d��Y"���Rj�i?AyyAB9����M
7�Ǜ�PVwt����I�����{�n��cG����Cދ�['���ƨ�Q��k�D�l�و�/�{��w�H��0q��3&�2�e�{�5Z�
VH��������^ɝ5��]y&����k���������+6@J�x����D�Q���@_w���O{���
�*�뤷�N������0��P(-�T�:�!H��&�ڜ�ؕ��["��e젆�?	���L�|�)�n��n�)j�'W��=��#?��	KƵ�����I%�5��z�1�v[�M��>y��^�<�6l�9Ԁj�?���KL���eXj��n_�L�_
w������/04�[V��VUji]7�{�1�G��� 5ȼ���Ϊ癨�F�����'��rD�f�o����1���7��7��5w��˔�+#aY۽�>U�uZ�*V�ݬ%�(�6D{��M����OT���م��Ι�y�͓U:�܀�!����+>��6�56�'���{�֛]!�
�Vc��!��3�,���'����(�^���R�Z���Sw�"tO��~�)�%����l�";�h����A�(}���ƞn�� p�i撉p��EK�i��c'��2��/�t�L]��G�D���F]�ðjr�:�5�R@#I"*�"�ῠ�yD�ɤ�����j��mDG7u*楓�&Z ���x;k�"��Eh�~2�y��0�~ ���I��6ߴ�����/���L{�Ї�N�ۡ�xr�{3���W!3V`��:���Gwh�2GxGȽqS�^��߮(�̻�c�L/ǧ< ;�rV��#��?����L`����{�x8}��	�/���URmݥ~X�q"B�;����%��Bx+E�n��콝
��z�J-�4hti�f��2y�*�8���I����/9��y��n�ӣ��G7o����)�:�nm�>P��M3��B6 �6~z�����n2lĹ���
��=X�q�FY����@P� �7'�Y&-���5�U�bZ8�Ѐlu6�� ���4��cO���28a��I�SD.��N綑}�QǪ�k�����)_�r݆��S��F�s�/!ށ���t�Lqg��0&mQ%T|�D��~m=.H��{���|ƈ���Y8 )���(���!;�,��Z�F��?}j�YeLء !��ǟ$�11a�<�n)(Iƃ������/��N3z"2u!�P��_p� �׶�I��G��j-fV_9|8?(\�������-�_:���f�Ԯ߱pp�-��ʹ��qn����u<wp�P�E⣲6���v`���gwF�jB�`]u�0�#H�_;�o��")$���H��fG���:�)���d\�d���''�_�pC}.p�7�!O�mkɛ��gK��u���K���q��C��N���Ҋ��ܿ6-_��6K�P�
듽�ËB���:��``���q��
v6��˪�W���_/��'��[�g���B����٬��}a�Ç`6��#�j
�x���UOo,&a�G�M���
;Uhx����_]s�EP���1!_f�=��p��nu���'L*�+�����P���3�KiN���Iv{���CF�Q�*��Fa�uձ�9��Q�#/�!�yV)�}�jC�.%�Sb��i�5�>����~%H-詗�>�˕�D�o*�l���:��K1��)Y���&�t�Q����yM��l�4�v�C�}s�C�*ڨߠ�S���B��C�wg���N�{��(�h�nN��e�*T�ny$��x�J{G�oܒj���'��%�Na��bA�v���0he�sr�l`(��
����y��ډ����6�+�~�`ߍŵ͋)��ʿ����mY��-h� j������Ȉkÿ��G`[�TCK���n0|P�e'�Cˀ�<.w�Jq�;�Rq�Z��c��7-�}�~��-G�4g�.��0�J��O�!#���R.)�q���y����ߊB}��&��@`P�t��!�y)%?^�y�y�~�!Z�����UQ��y�F(�kTS�&��eG�遀�5_�B��;���V�}�-*��`�������K��F�\�FM��֤����/4���k��qT��#� �҈��i��A��*9��h��^�hs��x���lo�J�R��i��9(<�1��WZm�M����p����~r�*�!"�a�ٸq��������o=>:'��А��	|8��W���vEԚ�Ǎv]�*%����D����G�H���żW7]�Iw�l;�	�e�|)4�W_�b^Ac�lt�M�����R�]�ݜt�nD���t� H�8+���}Ӎ������+J^��`��j�܆���*��ȉH*�"O���Ӽ}��j��i ����V�w^Wf��rʌ�C1��
�Pi�ڭ�yK�x��K��)U��
�d�
��}��A��ͧ���`Z(6Ԕ�0@��D�����j� �4�W�a����R��ү�~�h$�Y79�ɥ!|\��Cb�Hy��t�蕼�WyU��{c$~(/�7޵�u1
�b4�>� Zʤ���'�b���W������8�7f�	�z���Y��6��,є7W���6�'i1c$}HfSn��r�F��j?Q��62�1��W�);~�����趌.����{pj�ڴ���,��L��xE�$hC�k["�JH$�\вŅ�]��F ��
�����Q۴��:�3ljj����,���025]�w]i@Mz8K����2�x9�'u����WI���RT��e�Gn��˥��cc����1�-8
kZNZ�h���~9D����uu-m�|�բT�`��O�~+���PШ7y�F�$���.��7�x��w���[���}�X��tp�F�Ӓv�5�1������+޻�$D�Ԧ���%b4|e|�Z&�"X��i���0[.�:lC�>�k^ �4Mu�x�̓�ư袠)L�Ӊ��_c^&�;�P�:Y����E@��KH��^�RVqĬ���Yg**)�Ž��|�{�K���o>����0:95o��u�.kۧ�Eh���A\�Z��[(�8��Xm�����&���?*=b��tB���%#�n%�ϝ+��f����o�i>5q�i��ƪ�R�Ǻ 6W�|���& z$�@���rs>��zc�l=>Ԝ�{%�F;�;�m��Ro�cU��\��
�,�|�ނ��'�"!�Y*CÀ?Ml(��2X�֕�HhWՌs�I�	��f�H�Zn~_eg�������f�3ԃE���W�4h,}�M�S�$�ȽA��^���7s�j�Q>�@(�3jL��'�Fmgj��%�w��+8���#.X!��Ϣ�bP�{Za��qȚ_%x���s��������c�x��g���u�[�.���!;Y�eW'�����C�
9C�����[�$��[ݎ�c�#�E	�C�1΅}��� z�ұ/��{^�;� e���yv��t��M�7\4lS�gd7�{ͳv�n��1o���"��#�s%U������nt��g3��e���n�̀? ��"ƚK�"���A+�{��Ӻ�n�� x�Y�u��¯���Y������_T��ؓ/!E?������Ew�͓��$q
���Bs�r�n�M�*x�ZK˳D�U�-D���o�)r��"c	A�f#덛#����K/�:��@c����nAqEc�'}h0-p�{�5Nk%�M�kk=������Pn5Me�ey�S�C|��v�{��x�%��Rn7����yKy��/�������?x�(->J����6��EU�����Vu�V��R���Ds���R"�<b3?Ψl4\�|uxOm��J��j�ՃO���7�Aac6�[D3׽Zvw�=5�xuHM�9��cR��G�6l�<�v��*�ZN�ƴ���Z��j��Qu��*�k�a�ѽ3����<�X=�C�EQ�,ye6r�Z�V�~XLu/TYA9����h��/�D��_�F�>Z��=J�D��N�ѻ Q��ΈD�u���y_~��Ϸ��cֽs����g?��w�Zc����&�*t���3��(z�o��S���dp4�3U��8E����瀗>�'�$�iȚt�C�~B��N��f�P�x���`��p`��Ͷ�c�z841�Tf#��E���-[�A@k	�B�tYX��\��e��i�,��4��c>R���rvDw'���j
�Po]-��k3f�گ�$�\Q��k���V9@�ԛZ���x���n�BQ���-'�.����qV���B)��;�_�m0suڗ39o���a�ty�`�u��y�̳{�A�,yNz>>f�A��ab���?����Zg�$��=�s�o��n'�`_5����e���5D�P��kh��A���j7������D��H�3`;~l{X���K�XB��NX]�sxBs��A����<�Tw��\o���[���\�p�F	�
�]M�Δ�}/(�y��,@�����GB�]�#�I��V.��G3�Zj���U�!�:��G4gkt���/������~��>��Xb#`���p�����lV�y�uX���e�N��g3�f���O�������E���j�	{+��;e-��+m%_	���]�sO����\��9��\������9�t�lW��^�yIs5y�����\�8��D�G��F�!¦�Z��G���n�o�l�|�~P�D�r���m�#?_a]-����O��Y���_%���i^�:p��栘�v���t�:|�N0����)`���ϔ����C��rs�V��Yia-YƜ�=��n,��@E--��JM�K�۩������?��(��qwC��9n

�+�频�8(,vZYr�-R	���7q�n]�~�]�޿?[�-��6NT
�|������?i� J \V�]\yY8y	ޘ����@�r��}�w�/ ����M�<����F�o4}�A�y0�O�3u� �Sr䅴��g��ؽ�	f)IJ���Ks��n���5݈��<p�`��\������|�h�p��6����8��H�ubVVn�I����Ay��oh��	ݍ�;>��o��0_;�[
�S"�3F�l�.j}A/��0�������#&�á� �pcmK�i 3'�ⅅ
�6)�2�?�]��d)Y�~(��Ӏ�����%�������bmp��p����Qv����S��
֥X'#��D�s���L[E�`��dL���Q���9�X>�=��}]}#b&{&O��o^� �������Q�]�+z[r��T踢�u�?�Jind�Tf]��Z��b[蓻�z�[�,��!�V�5�*��|�����'����~\z�T�Щ!l���|���I�tHڛg�B?j̕��s�d��mͣ�'�[,��O?�Rǔ,3|�1����4�nlɘ5�!�#+�?�����O�g˴�W�'�	�}6C�e+��s!R��&zg��1G�{pw���:n��T��#��}�/4^@�56��Э���Pd^��9DوUNN.�_����E��~W�ӓߖт,t�DR��K��H_�4	!ۙx��쭉���yE/���J���ߝ��̟u�B|�v?�p��rt��f	���IB:�+X�g��۴ VƷp�bd��d������/��{Ȇ;�l����Pi�H�|��)��������+�EG2y��������I�-�1`��~g�r�8��10F�<���0�[�8��?X���uW<�b&[sˤ�O���bOy���M��|��a8O�v�����%�aY;p�� z7�^��R�rK���i��Lb]�K�iޘ����2�n\4�y�?s {�uqU����!��z�w<�Z���9�ls��.����c��̆SΦ��&�RW��'����	��4���zӰ��臼�*��7�^'���'l����q�ҟ	iǤ�(�A�@�6��\9�q�2%l�N"?����������+�s�'����H)�it۫�3�L�ה�u�R� �����2���Er�Z��$�V�f���Ɖ�f/��l)�D3�Ĵc��2h�|���U��M�v���iG'�s��g�v�S��j���-�r�(^!����:���X�'
?L*+`��k�ʹ��MV����O���Z����OY�G݅���	�&�z��X��H#ڥ,��y4�R����>5��K&gd�RP�a����c�M�����يo;��Ӧ%��R������?[4�BϪ���&~
�{�\����h��O�PG��JBώM�kXĥ_10�u��q�͎��D��nH�Xp�ķp�S����lr!�kEI��J�Rܪ"���"������sGI�"-��8W��[0B-�pHn�;����'  ��|�Ay�e6m��`�?�u�Ru��/�<q$�8�������9�4�<�'�lʇ�}q���z17?\J>W1�}�$\�¬��RN #±}�q�Hl1�g�D�꽯��Ҙg�r����i(Dr�l�J���wA���@^�I�ƹءy%��Ĥk�[o=>M-\�D{�3,K%�G6�v��^հV�j�)��왌~1����9��25|AZ�7��ئ<)�ē����8`���Q�R�?���f�Lɀ=�j�1�;A�MX��"�_�B��[-�qO�6kY,F��T�z4������R�iiCm�()22��鱠�3F#'�6C4ZMTJu*��zk�X�G���km��}�-63��0����U8�q#��m��t�A�א.Vn���99s�O�2©�;�?��K�x���~��Yk�k��s��.��ɣ���g����o�`�\�pe6n��Й@yv^-�q5��"�$���MǏCp	�񖛞?'s��y�싆s�#�R�1��T�v��
�^�X�9�����".�k=pڮ�ߢ��:�Sd�64f�9S���u7Xi �y��kF�	S#"
��&�8 (d��- ��T=�n	���m:�=�0��G ���J�g�\D1�R��dlt,w{}�#��V���7�h�ܠD-��h�SMqne�lr����# �`�R	(	��=��6���H�`��Ĥg�#3¸֎�&���D�
�撏��t�I8�5G	��*S`O���ݤ)8�[Ngn:��Y=�i��_2�oͽ;��{�0�ހke唫GCg�~�u\��r���=��o�;3�1Ϛ�������X�I@�Ԧj�$����a��f��f�t}W�\�7��$���tȫIl�W+�P6i��.y%�6Z@�a��8P}���J<��x!;�����*��������A$���ls����Ն��i<����^h�ٙ^3�x[5��px7}�@Sǣ����L�gi+�(����Q�6�B�8-�,��Tɹ&0��*m�E\پ$d�ͳ���C��5��V����%Q�gO�I,:>Q|�b@�*�3��.��a�"A���]&��>��A)Gۗ�O:��^����({���E��C���q��.���}�UD�F7�O?�廯�����F�S*���WT:br�;�O1���Kk����|�#��7V
���J��B���05Ȩ��I���1b
�إ�?*����������S�)�n4�U�j��,1ϓHM���6�诜9:�7�M��/mm7b`�ˠ*�V�����i�f��~E�`���� V{R�Z-ܞ^�1CbјLЩ<�t�W��M���R�r�!���s�	q�F�0��f���~�)������L$1�G����Q͆�h�0c���`�O{�RBfh���ic�"1���o!�ݵC�W���ީet�?jD5@�+�ͬV �/B(�Aw�{�ڞ����S������_F_&`�u�^n.̑L�<jXD�iK"�����oך�	���� �yS�Fz�Ϝ��E�$�S�&��&C[����N��)s���HM�K[�*e1�S�f�M]dTw�C�Xx�^p�9������k�]�M��n_`�Ѽ��6�c� ���sӮg�ѡ�
�k���ܨ���Y�љ'�Z�bF\ڭ�K$��nG�'�Y�f"�>�W� t�̧��V��Z����v!�n�ӳ��Ў����1�Ɯ�h}�No���ﾽX#�X��P�]�ڬ��^��֟�t�=g�kֆv H����4<6�ĵ:�ݤP@�@j�0xl7lo�lpw���R~�ڤ�R'<D70�pB�W�;+� ���չH�s7b���E���q�I��5���X�WY�}�I��:jv䜡Y���$	���5��f��ry�����ixW"i�l�-힕��q��u���+>�-��",.�GP3
�R{�>N�`���'������,|��.�Yʚ9���` ��I�$u3� �¹I�������2P����F�["�T��s���n�CԢ	�eA� ���f����=��~�a`��#�8�#�Hb�R���k�����~��xt�?/2J�����ehd;3�Suh� ����B���<��"�6��:%��I�Ӈ����0"��ߺ������~X?�l�4Xj���iv'�P�!މ�U#�j��7���i!�K�V7�s�b�Y�s�b����������j�ѓ����τ4/����O`/}l�L��U���� �c)�|يjaib��э����h��ޮ��/(�e��Qd���b<Lhµ={���y�,P겐�#�7��"��/�9�����}�Ufq����{̎.�	�;��7̊>b{YN?�8��Z_?��me��Z�6��}��Ǝ�M����V�	Y�񋓻���mc���Z5�=��.&�\aD�j��گg��q.NR�����t㸟 ���N��E��1�0iB���ך��}@�j�P���{��t����C��I�d�!5%��PT���hk f-�լQ@8�^���,Aáz��BdfpK^�Z��L�������^mWQ?����Î� �V�`��;C�K�::����[�~��p�w_��5IO��e���"O��B1n�Dα�6pA31L�m�5�K�}5h+pfh�"c2�Z��ӑ��0
��G�eZ�ý�E���j��>.�J��k�	 3@���*��U��: )�¢65<����P5��є���#)�]'&�$�&6��!���ӱ%�GC�_P�Ӟܢ�7�J붜�e����Ǳ0kތ�3���!_�AFaϩ����˘�06��Ұ��J�YxXL����|�D�}���Q��Q�R}a85Х��,C#&I��N nE�X��C&1Tv���e��m�{�Ώ?��Q�Y�j!���8�6r�77^����"�L��:�Ol���z��ٙ:従�-�n�VO"�F^���Ni�AJ�a)o˹s��3�~S�<����y5�h��>���°�ȋ��h�qUyU!�VR(�ϞV}�H�$=�t��5�+uZ�������L�Q<YX2����pxv`�ߏ�\*�bM��H�=
r��ҷY�0����%M.̚9� }��D��]����E6�:�q����\O,��]<=��e�P��g�&\��;�n��(~�����	����
��!!/��băKqQ�4��e?v���T�?{ֵ6��1��~��>u(2I���' �;èA��Mr�:U�K��$.�)�����U{��^8�u��Z��A�CL@��ݸ���4�^#��I-�ݼ������E������ �̼3��'_�gn���,cV�0 $?(�^i��߼�x������:A2�;6Dw���iʊ�����[F��4��������I��]�3��h�������W�`����¥���D���R��sh���L*�:��l�h�1¯�y�%�Hz���nPBk�m=�4Qk�/~����:CM-�S	ZԢ�'��n5h4>��j����^�n�p�O��7j�(g��>��Qv��\����愮�Os'��ky���P�F�=\0憐J�+k6M�Zk��s�ֶ��^�O�E�\�Z��y��aW��\���s>Yf�+�{��C[��.$lW*a���xe��O����˹-I�����B���4S��>��ۜ��$K��H���'�r5s9W�F�k���1�a�-�QY�
�w@Y7�NrD�ŁY�T�IEv�5��J��Es�t�g��cG�<�yu>��-no$�=���5m���H�d^�*�\�F{��R����<��l�%W�av��F�;��x *mI8�B`qJ����ܪ�g��8��|qt��(�C�Q�����>�3��U���Uo��l������|I��� ,�n,�M{�S����_O�\�p���0��c�� ��u²�XT5��;x����EB�����3��q�Wr]�V{q�@�����k��>�߼6�O�Z�v7H��܍]E��p�R�pm�U���J��Y�sł�lP��L��?9���܏��m-GtrӃ�}�L�7�?}՟��yĳ�!^K�E��A��ҳ�B�d3�"5�?�~��䳓q��ǚ����s����Ni�
}\B)*+��1���I�!R��b'���Ǭ*y�6���2��u�_*���N�l���$]m��� �K,�C������z�<�WRd�����F��q�z��M�Z�;�s`�� �h�qo[*k^�)6��w��*p�*��M��� ƭ���θ5ƄZd`�HE�a��B1$r��&d�lNFx([�P��m^	�����s5t���XN��,�� ��h7�E����Α�Bx��@�������N�=v��c����|�K<hϒ�R��͕7j�r)T�< | Z۱��4Ȑ
��>)��p�pE��^�U[�_D��9T���
eD{%\Y����$�zѥg�� l�Q��3�����q��rPJ��������hr�P�^X'1�y<�"�v�-���R �����J����ť��q�b}�xЯ�튛~'�}�w8��MO��Qc�ǽvAuQ���s��� �ȃ���H~Ȥ4sձ!�<=Es~lM��𺴕����	H�r�&&�
0S�����+���Dx����&ݻ���_&��PQHި2��F�)����ͅ��a[��	��MI1��Csj�m��KO�-��N��$�?1����~>7�K�;W��!�+���$~�����\O�ͅڡ��"�j�	]��_�inɊ;��ki�y�M�po>�qI���N��fq6������:ޜ�)�NQ���ؿS��n؍��]�+z��⹩�w��P"�տ�:6�ۃ����P���gXkg�S)ь�覗��⁑���뉝M�h���xV��Ĭm��ܮw[#C͝����ƞj�b�����*N�e�6N �h�H�yG�����_�!��N��!���Q�w�=����·�(���1@�0�q/4՚���!ok�z�����ً�S �x�7R�|[����D���t�gSJ�m���m[uŽ�9Z�U<�8
)�r�|������"�@�J��EnW��,۲ں)>W��l��l��{�y��K39z�c�=��<J2u����_O�Q���G���0�t1]������W���x��b���|wĆU��k��0Ԉ���Aռ7|5���D6g�����Z���\5���SZ�!�&�+�B͸D�oF/>׾��Ul-�W���N�=��T{M:�7��ςJ՝+n����v�sa�/��h4u0�kr��>�V:u�gew2��iZ�r��ɡ�*�o�Ȫ���p��Uq�6��^�O�zS[�/֕���X3��1w�o=��s+x�ݪ�����!�_4/���)��^�]�����]t�������U�n=Rz��94�Y[/P@��p�\ �vϩ������+Ԗ5�� �]2/���9����K� y��HiaAX^�W͗Ww����񾵫�>+Gq5����oͱ�h�6CZ�°��P|;}��1��7�.����u�)H�xp{�����X����|J��f��0��
r${p���~���hCk�i Ezz|6������Du(ո6���zU�2�4og���8�ސ�E�JgF,x��X��l��/1ꢍvc��:#���)'�7�D�]�k��mE�(��N��K��G5��a���ԧ���b�\�zմ�����Yƍ��M\���]x[�쥽�16'o@�y�_���K���2>�>aea͟x�^|b���k��O�u������HE
d�@]W�c_���ǒ����A�gM�'}K�B��Af+y�����T
�^�FBI3ߟ7Dt�=�#�vYΩ�f�O�'v_;�s;��
HD�܊:u�0��U^�}} O�
&�
H��pTY�zA�9�{w_p�%�&�Y����?�Y� h�*�����7ay�{K.���Y���d���uu������9��|=����@. �E�q����=0B �����V��|�]ɂF�E�� �?�k�{4���`j�do���7�' ����*z)�p�S"���^����]+��a-e���`0#+���<�A���v��(��^��-�~"�b�fF�݆X|��4^+��P�B@��n?H-�č�}���8�h�^3{s&�\��i"U7��;1�^�s?m�h<��_X���?݇�����5Fz
"�]�&K #5d �B���l�r�nϫQ[���>f!���d)�Ve�W�%P�W�����Ѵ'T/�Z�Jw����,y�}rթ�J���`��F���כ5�`_����nMI��\�s���PK   ��X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   �sX�@M��  2�  /   images/959826c8-9748-429e-bc6c-0234da684cdf.png�y8�o�7|[�H�"di����Ki��-ɾe�)E�%d/bb�%����c�Qvb�c�����<���{�<|GG�q���������u^t����� A�ʵ+���h��w�'<L��{��q� =%���׊� (gP��%M��߽�����I�f�rͨ�����6G�0.��3��g_P8v��l�����+��8���O�':�ٳL#��/Kc_��\�U���wu~�4�@{\�{c�
��=j<]����˯�U;vj܃H�d�k��ghe���,�UJ������/84��!���Ϳ�˂���xiSSӊUL�G�����4q��w�ou4����7�:V���So������!u�ݻa�^�n��I�Oed��A���h�5�P`��[uG6������7بݠя�Ү����d�2��W~mcy��ˣ�a}�%DE����"+���G�'vmu�<Ƞ!���O:�G�'r����P[�<f��ׁ�'����Ms�V��iE0�?G��!��|�P7O&+]�:���h�K|DC�.��Z�,#z|{��#���u�E�O��Ĵ�H��WU�+����n�/Xo�pgC�J�8K$���b��m��
Y61X��e�_�ɫM���J�����S�>\؄=�~�޽ӏG���͉��D�t"!񕄮,+��E���h?�����"�w�ޚ�x�#�b�H��h�u ����u�K,�%��c�4�_Uuכ��Hӌ,o�f���:�T�[�����b�1~�G�/�ǟ>}b�7�e�w�Q�j�F�wO�x�ެ�_����u��d}�gL)�,XPY�R�K���<�h�)O�-��c����S$j��pHV�0'��"��}d�m��n6M���^�N�v�poi�c��m���\���Ϻ��u���Kh�{�\Y��B�����֥�~�q������K�y{���l9׶�?~|ȥ����(��얰�����}b�}����X<<��zm卑��;ʉj���S�I�@�3,X,���̳{I��O�un���Ȫ�EG�<'XK΅��Tr��j��f�}���6T3l�\��I}k��~Z@y��.����;S�PM}@;߯� �lH�IvBؖV,���1x�y�FR��ԁ�t�A<~x���.k`�̱��l�P�]k���+S��e��ꎿ�?�Bl3%a���/����=�H�i��O,H��V��z`����%�� `��`�%>V�ANZ���i�51��.=4Uvv�::E����?FXS���ZX����99] Z�OI�=w�-��}y�����ə��Hq���bȡ�<Y��>�U���*<��q�Ϯ9���o5aެ����8�@�x]�K+ 	��%#�`����iy��y�B�o��R���'�X�y��d���$���v�Tݛ?ћ��=�xps��g���ʐ�w�1�\Q�呣w*H��j��g��d\���9���t7�����J�/���{���L�G[��bL���3��27��x�v�}G룆�\�/p���Ő1������ N�#���f� ���Y#�$� �˒t�S�s��LX:���,�(�5��OHl�c�u��;��������GF�y��G;�]��x�bf�}�bځ����g%Lnn��s��ߨH<�@p<��%^���΀������^�~L��v�U���y566�M�	����G���qX�� P�j'�9�v��6�W���Ivy%��,7����aڟK�l��X�(H�Y*��L��1�S���CP�8D<}�`��|k����A+ڴ���T��Փ�6Ω�b��>�Lק�����V�K{�̐����RܫнHc��K]]�xtJ��;�,���4p���#K�+�����W�O��|1k=Ǚ(�Z+�f�x��)))�XHĆ�a�w���t�^s񈏒J[����0Jl���\��{+�\��Y�[A�+��8Ų�J6ES�j`sK�ðڗ/_L����v�`��OgɊ�c�i�s����[���ߘ�##�����RZ�X�����c����������Ą4�~���2�{qq�E
6YYJL��Hl��`L�pp���w�ڦ�J��ϱ8�SM�5^ͮ�G٣�.��u��0�X(����ٴ>��:�Y��)���EH�����>k3uh�UYx�a��I*^�=����(š��������ރ�>>>�
��Պg�E�Y� .ZI�N��\B�}�p'ҿVMIb���j�]�!��9+ǵcb!K~y0��b���:��o���fQ�nn7펲�\�e��c�l������������3a�+���s�%e�9,j�ֱD{{�'{��5Үē$���<K�#�;�eH�vwrr��_�Ԕ�⯽.�F5eU�(���H=v����e�Lo%���k�����/8�<�%�����[�s8�WR^m#���R4T��&u�	�����xx�
OW.Wlt���'o���󣛾k��}�n����>�m�Ԑ�4�&�k	�Hi��*2�_���1I�s��D:�L�N6�Yc���5VRW8���Ȫ�������N�sl^ ��Fc&������z�q���g��	��4nw�$���sMiU2:��z8)��$��D���;����y�Z�zlr��mps1��
j�Y���#���4�Y۾.e�{D詁�I�Z���H��GH�������ĢJ�e~�)��c-����)��7攔F..F�� ���$�Of_7=_5�,� �ߢ�r��iI�W/�������n �R_/^�7������o�8���<�.���RF��W>	�>�x�=�(_����E��O��M�pMs��/s����N��0�1�vDBJ*�._�5/�|���ي/�U�I^��HkOsKKCM͕��{��{O��/w*$nR��d�ͦ	���A�n"���t�$��>OTߺ�5'�[�lI����&b[L�F�A�<�ҧO����K����%�ɱ z6[��8�y�Q�V��`�f1raK4ɏJ�8�DwQ����Uz_�Dvk�Dh�.s�Hd��|^�Hx����(��!*��/_:����GP�ٷ��b[���!B6�E!&''�E]�v��}� ��I�DD�ڎ�S��?FGGp�t�te>nС�q� ?�8g�&�k4c��p��#��F,��EN��;=HW�>q��������K�����Q���Z�X��]�e;ƌ�y�z6��y��Zx1	L�)��j�>�����ז8�npkgV��	,�m���Z����I�"`�TD2!6=@�A(��v�n��ZZ�O^p"�\U\�P���@��[}��[\�|¨��e�u���=3�Т��XZ?�0�����[e�f�ܮ5�,�y{��ي �Vvs`����k:&ff;��F I�����LD������?~�uf�b���?��֦]�����w�`������Z�N�S�V�v��y�wA�Ǒ� W}o��H�L�PA�Qcc�<V�|�`,�}��y?]�b(
�W����N�مL���略E��ظV���n` ��Պ��5e��;�Ji�s��4Q������������O�����B<:�+Hao����@���hg���z�d����A�#�@�N]	��� �.�9�<t,���(��I��F������A�Lٙ���#��n��x�~G������/��s056���r>��2�;d��K�SE����s��CYIR�S�wOq�YAv�j��ާ^��D�4�)rs�Y���L���R�i�o�ؘ�lB���VK�*���(5�;,gb�v����$���떺�H�}n�{gL�v�Jp��PR��!g�O2s����` .}��!؄�4S��i��*X�!�=s_�=��W���� >����ֺt��_K�%��h���~�5\Ʒ=�ЀΩ��l��脄ȴ��9�!��3tVx�~q���;���C�Fک���{������ i�cɝՂDjȡ+(�5�]i � g"��K���nF�>Ȭ���Xk^tČ�8'Ѿ{c�c��ĜhF�`��7	w�ݿI�{.�"�R����A`ҶAG����8��g���&���5I%;V2���[�291��S���ɬ/��Zeڷ����kڕ�8�E��)�J!�H���zʫ�|�`�m/��U&���[������La��U�օ�>�i��8Aߞ�<�(�l�׋��I���BCB�So��B�Q�&I~�7��}Z���1�Pj?V�p��V�* {���`�n:�c"��s��n=����&1��~Z23�[6,L�X@���JFFF� *H��V���@#/^�x�3�(�<F��9sR�gy���p�O3�s�hR0l��Ҥ����뢓���]~�ctf0�xק�555��V�c/��N�홲�&2� +��g�{x�<��s)�v5�U��^�{o[���ii.���V��i� �q7��"�AU��t�A��� [�G!	���'�z߿�l$~}�2����?{�[{V�W!���I�(�"�� /���<��d�������V�}�����t�~2ٍ������ܜ_|��w%���{��D�(�K|ͦ���4m#��ͪG��|��C�B~���Ƞ�=u���)xy�N�u�Kf��p����f�V��oF$U�G
�(hj��BV�Y�W.Vԁ�l�#S���&cC��Q��oe8�x��*�������y��I###��El��	�勥7��׎�w��S�`bb����8�Է�\��l��"�Z�	����ݓ_�|@Hu���j�(~�~z��I��)|~��@�q�~�MzUr�>�-;TG	J�=��o�&��$%
�#W�����7sss�b�]���݁�� ���fJ*6`j``��t�i!�R�M%����]�yy�l"�������nڧ��m&~�њ���Z��-�����-4�Ikv�����;(�����z�(3U��6���A�@Dn�3/K5���߹���Ձ��\9S+,���	C�,�=ǽ�}�r�Vtpy$1lJ �EA�*!ː�W��,5$R���S���z�
�[F��������z�x֓�FTގ��$/e��^�w�����̒qA���&F~��`�iy�gs��5�l5��M����.�R��C�I�	la��(dD�[uݗ?�{�J�+�)��ӯ���Ӗq�
ٿ"�����ˣc�y��5$�����ﳂOl���;�7��K��]���Z��L���S�����ח�F�EC�m�f���C
���񊊊SO\k?���p,a�n��W����p}��{�+(��Ⱦ�r}��!�rm��I�]�!e\;�4�*��aC]����ÄӤu����ULMMzlY�Qq�фn�����`�ɳ�2+}�s������--��q�=8FG���D�m,�E�.,6��ܖ���2�)���'�9�k캡��o]�܇Ji�	j��s�*��D��{���ߟ_<�{θy;�gǲd�.d�R�\��nƍO�>7GuA�y��V��b���4������������i��)A�f�����bוui0�D3�)�:O���V�c������˯v���S^���R��	�޽;
�W����xuy�nC�D��|+{=�p�X���9GG�Y
��жbٔ�/?I�Goۘe�h������x�H]~�})e �J�Fl�W]�_�WG�Z�|/�[�4i��N\�(�Dǫ7�(����!`���a���ȕ��C&�35��r�H�Xb�:��!�V.�>�f��h�O��F�|b�Oj(�mZ�2�J,���'��K}�Q	D�	����-��Ve�������أ��٨檱H���e�<��˵���Q��������G�
 �\z���v&�v0M+W�L�۠�t�5��=~v/9����x�ƍ3+s��Nx�ʜ1�6c�2���׻�Y-`�P=6%`W�3 ���w_���a�u��zwj7���������I)�>zZ]F���硍c�~t�W�.6a1���ዓY ׃7Z~8�}9�ĵ�8O��j<�TE9�g��X��t]���MIV����}Kŋ?���S��l�]�+��/˫tؙ�׃,O(�ȸ��;�4�|@����6¥�WI�VV��9B���H�[<
����m�E�������[�����<��l٪έX�2��M�'n|��8Z�2�;0he�ڝ�)�g��PI�(e0X�b	|�XXy��ץ'��
��3ÂZ�d������)�P� ��>�-=�^�\L�]�/\yk�}kk����'��b_afSU���Uc��w���Y��Y���SK��Rd�����L�h�s׃�� ��3�,�U].�]-Ԧ�!���8�Y�%l�Ĺ����e(��6���1��l�B�dB�I�CE��`�W��b��N<����p��Tk2�,��{=6�$o�g��������}�C����y�����APra���w��YM�U����[��U�},Rr���9�@��ZldL�2Bz͵�����Nא�}6Yq����e�/� -\wJn/�������h��ĕ$)��|Refb��ా<�lW�9�T����`��b'x��}elLu^DvH�4��HՓ�����B]Y�����ò�~��?�z����O�o�d�'�d��(�R"q��AxG�d�#e����U.��i�r�j�_D����,!Sh�6cB�����Ǯ��+4ؓ"���kVsIY 0��}�g��=T�6�7�&��ey�@c��t�*2�����d�0����P�>�ȶ�)�Wa����S{S�,��_��a�?X�Ļ�����O�M�k㊑�\�yf3A�I���仱:$d���W2km�4�U?����c
7I�,����
���F�X~M�,�=��{M�ϯ.��_�W�b.<٘	�&n���j�X@O�88^�K�J����o��'���av��\A.��s1�6��'�s��Qe�jO��K23ղ�+Io5���Hhoui��W�%���j��m)Q��+�~��]3��F�-�����vo���E��mo��T^�0����R_s�U�.�̘���.j{4���9�J�$�O��U=j��|���=����&&��Ls�qzo]������ole�Z�ck��/g�����8�g�H՘�W��E�X���G9\*$���Mb�o;���g5!?����x@�(�Ñ	����L<���4���p���ㄡ���j������g�p���t������#=��g������e?w#��Ka�y�5'���WN��4w��32PL;�֫n���|ã���KҴz�0e�E�IH��ڠqa�^�P�$K�}-���^;q Qm�ʧ4�G&����p�ƽ{�~�	�����Ync��Zs2��c���LoK=M�M�<��k��ﱚ�L���tL�s�S=���Ǖ0��G�����C���0���u��j�዆~��.J
�Z��ү~��QƧ��,�w>�P�+�]��H~cm�u�W���݂�S��zK����*a�ONu�����ui������'�e6^N+���z��d#~���1��^�}nf`v�~݉�{��i�ML�Q�L��ӗ]��Jr��}pP�Dֶ�׭.E1BP̾�:�Cvə���`��w�j�t���n~�����%��i��dTOx��:�V�k���XE�3f�W�U�Xm�I�uNZ�޽�C���V�	��6R�F�ʂ�V�0?� �+ԠQ5e!#�sڠ܀�3�4un����S��@�a��-�w��Q4Bu6��˧!\wD�{�T'̾)F��~�P�ǖ�j��)��)��dg�5�
�+��<SP�g���尟J���%^Z�c������5_'bo,��@#CW��|��'1ʌ������@H5��p��4rxF�^$H��T^S���D��ҥ��W&�M�a���[\��]55%.w�ܗ��,?�أ�؞�u�v��v�wi`�'��1��&)*0i�ʳ�t���	������x������ܧ��-lm�D���^�<t'�S�0��q�J��l"�С��!٧�@�B��i��^um���|^԰t&���n:�߿���Ʋ���q���܌ׇWן��a��b��Ģ����>NY�_i����J8BG�����O�r�ј�/�i,�jxX�쵅�޾L`��PXn���K,^_�|~��xD�-[c���Ox�)����+�>�Ś�^���]�"^���}��5�� �Y߾�U����� V�jh==~�[�DCNK;-�H�&�C�?W�g�:�Ww�+�~]�%k�XEKll�����LK��]ŉ�a��Yd��_��O�JH���:%��'p��մ�@r%�v}¥��P)"U�&�|�/��Q���ø�:�������ZQe�����ӑf����訇�랏��n!�[����Լ���GZ��?̦����' ��
�Y��νZ�s+7k	 ��K(���b��&d���V3�N_<�Y2c�4cKe�kv�b9ܟn�y����sÍ�Do��ʖ¬
]���Ҭ#��XR�n�������iu��'k��k��������]��P*~�s��<��T�9a�i����w���T2lZY�}��Gqs�,4sL��P���#�<7�KO�� \\��Kcm�������D���j�:��^?�5T���~*�1N��Mş|]�\����m�B�">[׏~+tP�~10�����ݫ�p|x��G�y��N9�i��ӵ.88=L�X}Z���\e�M욵�Ϋ�) ��$$�����{ս�H�%ֿ<����ңA�V:*��|)y��$��c������y�.��ERT�{|�(�����j�~����L�܏?�7�c����*k�|�~|����E֬,|�uFr]Ϸ\�マ���WO ��9s#f�lb�?H�����n��9���A�p��E�����ʩ����@<�'�o�W�M�RT�F&^z��N�T��~��O�K!x�~L�M]��x঳φ���~��w_�j������
9K�k���0'�3*�Q��`��p9It�@Q$7\`G�h�1mM$�r5q�'s˜�A�zp�9�M�b�]i�r]��R�Q��;���}�aF�UK=Kӷ��LgaQW�C)�򓳔A��`J�|=Z7�!��d=`��Um!(��v�<[%+��t�f�w�Na����WeE�E}'�Y�W}ks�&�J6=T?���+�U%�[b��EC_|�'\���r��< ��T\�j�!�\�"QOEjrl�bߣ�RT������I ��QG�ˎ� �H�.�u>��/����1�Y:�x<����3��\v��r��4��"/̷�@�Kʟ��璴}�[ꪌ'��.^�ny�>6λ��}���SQ���:��TG�.��I���=������d��K��7�J&���ȕ�c�����N�+���BϾ��a�T�GZo��n��
��e�܇�����>XP1�Th�WB�+S3�
-=F��F���<�}Ƌ<�8d��$�;�� \�}��Tԃ��3�L�WX�F�߹۸��j&tvv�|��^�Ƶ2��t�@r����g�V6����,X[oMvhՈ��W���{V��H�N�>��M��n�vT�2�H��z�A�x�AhO���?�&�-�ŧv0˃k��s oB�ƭ�Y[�gk�%w������f�12��	-:	�1	o���ݡ��Tb���� ����b<������a2�� rk`q���Z ����a�T�éOQ�)��x񚝍M�I�h�F���<�q�fϧ6n	I{��%�ߊ������ɂ#��^3W?��=Aw4û��FC'��5�ܤ(S�����m�2Dz��u�?�)�e�zx|`���g�#���$i}%/�
�WI]r��t̾M��	��N!�s/����񉉹��&b����>cs��4O�63L���gq�3��~�<;$
wF��6o@���{]���'r�����}CR���/��Y

sR9��KV�d�z����"�p�P�HDK��'Y��H�ƭ�b4������s����[J�)�9M�D�?y�c���,��7�t|�:v��O$�����b|���n�gu`��Q	��b��4Z9�f!�@s�Ҋh�X��Z�q/c���xo,��K]L����*��~�w�����T@�.Ү�-�du%#֣�q�F�o�6����H����-����sL8B5!�$��93�9u!K%ޅ��!����ϯ����?�ʱ����[��'��#Ezm�;7���vp}�Ϡc�y�'f�9V���p�ḫ�7�*=�lNm(mi�Q����6Oi�z��O.�m�iT�*[ed��1�Y��w�p��}2�ߒz�Ӊ��P�a��}�Hz���@�8`kkR�}���/B����M�'#+JΒ	%LAe!^����샴ӑ@�Ŧ���W�9�?��b�J�p��_�R�����p݆�ۨ��̓�(~�Z���B7�>ĥ�0���]:��n�{����ٱ���I��E�?��>z���lg��L9r$��͊�d��Vq�&�f�K��*Aa.�2�2��
���[r�������>����٨�E��)����0�ơ�ڧ�auڵ�9+z��C{QT^a\<<rY��D;�y;60$�X�*���!b�F���M�P-W��U�����>��o��%$�~��[̘vK�ya�=A��?<I�=�5��E�j���Ɯ�G�Y����w0�����䢋������x�����f�БdIS�3A+@��Rڴ^�<�`N�k�8t��v"o�WK��aA�c�,��Τ��~E�����z��j��! ����������1�|4�SD5]�v���m!�n���{��*�P������?J�0�]FFF���{�������S0��G��o�_��贲�r@Wz@�;�c�<a�G��
/XP�66Ff�Ú~�-��5��vsJ�L�X��;���T|G�UĮ/mm|�
�:؜x��G9��g2��y�~8���ҫ�E<5��
|ܕ�)M�'�6I[0"��N�E�T7h����oq��u�~H��;�}�X��gx�$���j�h5%.,�8#P-/BB������J����[�,⑀��;Ԑ�3d�<��c�Ζ�}E*EvQK|��*¬=�Zj�k�=�Yj5�����[��U�/I�%���M3���wI��q�ԅ5��=}�~~@bF&+�'�l#$e*�^�]dɞ�G���H� �;�$�@�x�
����ٚ�S�2ngc�wY��Y	���q�9M�uV\k�]���l�t�h�1�-b��I� ��O�e�ӟa�nO�z�Ɠ_�M���Sҕ�!�r�#��4����q�%����%��j��T�ii�M��	��'�%$�U�N�L�O�|5椫����E��ˋ$;�.�D|������M���ˏ����1Qݳid�Ш[�{�d�u:�Q%
��\�*dfM���1�z��ߕM?�"8~�!�����>�9���80�����lUy�ؘc���oi�Qڧ����B Aj޺�� �<_�a���?�^L�Tl�\���Y����(�K��)I$Kï��_[)	X���`�ّ߿�*���m��}��C���w�b=��૮�1Jp����*��Cg+� �T�P�l��>.ƃ��%�.����]���7I��a�����ؿ��37}7�;���
H�|�����z�}S���2��8���W��c��洹44B,U��_�^����� P����b����[�	'�z� c��x
��H,�V��R���5���+��wQ� 9�U����}`�P9���Z�i�p�	g&�8^��)h�'B#�ԋ�Z�+�x�� D���*T֗!�H�%A�ǥMO'D�Ơ8���z�q}�M�3>tR��d���vV�V��j�(d}�e�d�Z��=�|�f|ֆ�A���{~�}�����@l�C��R�G�s�i�0j�_U��H��d�x����
v5N�..�9  ]A�mC>����l ����ۤ�Z�ѕ��ڡ�|5�x�x�s/}*��7CaiL�x̛_H;`�u���Z��3����P�h�������/�<�5v�v�����dL ]��
h���+Ԯ�1��fE���� fm����]evw�}4�zoү��*a"TO�x�xW��l�7MS0.��f�ڀ�z��c¢�̱�g�Z%��*��ޠ+I�DbbːrDzs�r�&�P���!�����5\�v2���q�p-���	!'CQl\��q����IUWi������v��3[G���fe��9u�MD�e�g����g���80�_���tP�MOO�O���]�;N�&��XS}f����\��f��4�v�J��rr�P\J)w��nDw��+��G��&<���zW�<d)�|��)��+髧ix��f�S?W����� ��j�����jp���h5�"o/{�Je/��4��;���>X!p`��h7�®c���D+�>��U��5 [��=���7C��h<����E[SS����=n����h��Y�v�;B����ǿW3�[��6&mװ"��#�۾R�Cx��zo�8���!�lY?}��^�^hr^^�����R����
?U�Μd�h5�/q�/��n�r �F�2q"�1�?��cW@ +7˽C�ob�mgdH��w�P��6/��#�D�|�ؕۤ?�\�M��h��ߍ���R(��s2L}��^}��-�q��Q.�g�bR�Sy���� ���~:��^r4�ۍ��+5~Ǐi�թ�VN����/~��j��	���/���4g����"|�,����ڴ8���n�guq�?6�����Pl���"��+Q�I�~�^��A�E�6ϕ�5��o7�z��e��l�ף:��S}�:R5%�!���u-�z����N1!0�h`r8����?5^Q�����ԣ\������J�z��xC�0� E��߿3��%C�@vӺu8�����T�˾��k�BnվT!�0n)?��9��K���zHX_��a;����*��۽{�U��"�{����Y���^~�bS�
r/Y��Պ�:���*�?B����N��b����t�Wy�
R<��}��� ���5tt���Y;�I��tl�T�/˭R�|�˱�:X�IQ}�t��d�ӧ�z�4����&)c��J����[K��b�Ch�����~��H_�)�\vc�D.�BIs��XP�K�Y���3ͥ6z�u�H���|uuY	����9|��h���
r33�Z��%��v�*]<0o@L�͚nmC����j�4���F���*�I���f	��ق?����8��{�ȏ����Cn��{C��Y�Ə9�v�y;E<F�O` �6�ƍH&�÷��w��AnW�e�nP�|ޟbZ����b
QNg���Jئvn���_JѨv(��*�(�. ��5��ojL��pa>��~1�q��ߋ�����G$tAB�J�h�Gp�F��&�~�<�7}w|/��Z�f&�e� ��2�)20V��iOs�o��wpJ�*�;�����R=�(���&�ݓ,���t~w"��*[��%�vZQQ��h[(oe0J��dTV��������G����u[�fꗪ���w�O:����0a���v,���KC4
s�@� C�)��Q�N'Vo�V&5�G���w���|�������\;Z�@u��k��Mcu͟P[����S������pᇿm_�}�!���iȣ�kZ��w�E���Mc���J���q�}�f�
��������Jf��ع�8��^��A�����9iq{+�4��F����l�K��� Uޯ]79��Ḣ�3�Y|(+ �w��6�f��u''~���t�/�ݲ����_ׂ��Pr~��~d�V4�B��l ]���ֆ��D5n|*˖��9�}���j��p#��饉�������'�L(g���.�0��~::�,@�Wep�?W%��D@�7VB�?@��S*��7n	�ӎ*ۓ�5Ҝ�t�X��������2�H��2B_�Y��)�SC�ɱ��?����eڻW��iP`ŗX�,�I\OѸ5��}�֯��P��e˻n���$�H�ʳ"�#~J�t�1�> ,9��F�t�����(�s!�Wh�U�[�F+�~9((:�#:..��Ai+���8�^ �js��_.)
�P�Ɖ9��ޛ�Zb���v1��K��>�]#{��0� �/w�RMAnɺ���%j[|�y��N�����Z}�m(�����m@AȌ��?�h.���u k�����A��S���n�{��#蝻5�=�1���[��E�T���qT��!��v�g6�� ?�y�'���ύ�o��ǝ�n5�P׉T$��X��y�L��v>nyy����;�TMA��������`���Ӧ1���No=�3�"�˺�W�@.��G߿}�w��//o�q���ڙHUL[	6>�܁�>b ���Wm�D�a3$X͍#s E���K7�Y�����Ի���U���^_�8�y��]^O�Wk��NA[XX����}�`R3
��=�N�:�[��&�����ML�����ѝ	����b/�g���>4[ �};2�(�,���?b�+�P���
��Ǿ�xG@$�C�v|�&11LЬ{��3sGU�?�A8�9(I궃|�_�亜����/o��HzpwjH��Έ�I�g�-��>8�P�d��D��[b{���~_"��C��@�:'k�����`rٖ;��G����B��K�Ɉ2��w�옝��1�;<	�N�H���y+TԶ�u۟8x����95T�g��1 O�'��T��ظV�䏺+O�>�&�>���Y�s��~��w����G�>~�� �3;ʹ�y��X�_a4���&�
�\�1�shn�|��I���
F�AT��Rxa1�������y��P]�%�����/�\��rJrH�H���=�����ii�<\i�A�-xGP�&��"��훦���)d�ó=���n�!�����!��[�֍�.-5�p��[��U��d�F�wF݇��UTUl;�B�BPh4�6��C��׆뀫|��ԙ7��w�&���a�6��&�$')c1 �"�m}TQ�#��PO8ؓ������ u������u<�~]A,�w7�q(V�	�G&�_���C��%��A�'�*bJu��6�B~BX欼����]ʬ���]�D������[���&��jz�N���;�6R��Z��*e�n���/��ǵ�|W��*��Y뵴ҥn����.[�Wb;|7��T���t^�ء:���5��r�~nt�-uP�I�ۯ�菞x�M.Q_�s���t5N��E�V�h�{@�%�V�n��$u[^K[����Mo�%C�B�F��t%�3/.h����J��R�8����|�8�����J����3CR�a�ҝ�Y0��_�D���t[(k�J�����L�Ȼ(�l���w�U��<k [�S��]�4ӛ��b��,��t���/8i����S?��ڳi��&+�c��|`3�|�ji���.��v��<����j��	����ͣXMC��7��6�X(�B�wf9j�R10a��!�缵]��&��!yZ��j�zl>t2�s�X��H:��O!8�6:�%���P% S�^�L�?qq�\���v_v�df��F�pI�`ie/��ΘA�n��Sa�%f��5�zz��}.���W��|?J#f����9�|����(1Ӄ��V�Q��y���+��V�C:�ĭqî\�pj��p���2�t@2�8���$q.��8^]^�hX�ѧ��W�F�����]�-�θ�k����z����Y��4�~C����)��ު�-\�G�F��r�AȦW@���[�G̈́����X�8Χѷ%�4��d��m�p	���=!���^�^�,�oE(X��_V7	���2-9v*�����{�o'�㨾�¹�[Ӽ�a�e;��?�}������
<���:��>��ޯ�:,�8�D� ��b��u»;�b��W,�;u?״Y^�wB.Nnu�Q���l^�ZA�33mҹ���C�k��ZA���֝��xȷ�{�߃�����_���!q�Ǯһ�'ۘt5���S���]�� �4|	�j�*� �>õ����8?h����Be�b��Vp��eg��Y��_��3�R929T*�:��	�c)db�$C�T��:\����R�g�r�m�/ɋ�0�,	S���g�K����aÊ2�������*?)֪B���;C�$w��@x	��x��%�R̋W�J��P��H�v�{]����>�?v���͵%R~�56K�������o��W�K矐�Wg� e�t��m��Ʌz��������]:����x*�;L~�LiU�Q���C���6�c�L�o����6���� ���#>_8��}�Y��ȡ��ag���T~%,U��Qz�E��`�xT?��,�-�v��Y�x�MZ��5��T�	�M��+@��y�]6���Ҿ��[1�6���ݽX���x�:,G�.��x ��P�Sn�9����Yt�>�`�yăW���|XO���.�����o��g�b�1��,wm��y�|�C_�Xj,�ʋ'K�۴-����l��񭝫xJ����t��v"�g;��G���DE����Z�0K����"���� A�=��_�zWT���o�u`�jC~?��_��=����{�߃���� �MK��i"w�ʝ����ɷԺS���N���8�0mzs˥י�q(�n䙂Τ�8D�Z�6ð�"�Nn�����'�rv�y��-5n��XQ6Oʸ�x�WM��<Z����
�[ا�໾\�x���(d�3{=��k�k(�s��&�2�Ѥ��Q�!Lk����o����`(���C��KW��ޏ>.�Z��X���W(��~3��;�]f��ϲ�?�`���	ʚ���>������`�Z=xD�4YN�+UK���{S��=ie(���n֕}O��3�幑��5��|�:�2�����F�J=��g���a�(��~fU�I$ ��]��r|�e�t�()�o�d��e�|m���ú��s�m�rNi�����fR���WH��b�����Bf��(�Y��C�[�z�N�}~�%�.Rj��G��6A�RY�Ae�N��¥� .�S�M�什~�?pa��&�7�I�̥;ϻ�l��d���]��/vc�K'�3W��~7	CJO^8�[�ላ(%U�z-7�Z�Q���9^Ct�����Y�:�Js%���܌O�\��v�s����Åǩ�/V���Syq���d<�yN��[�_OfЪ�*s���vU������(�µ[��S��~E�!~�ɒt�����:^�2A�gbL\W�VZw}�������3������]
��7&`sO�Q"E��o	��Fh�yO�m��k ��D�J�����<�+��rK�����+���$3�M�Q��w۶l�K6 c�H,��+9gk�Q1��v�(�M4d�᯷�p�>'���P��Z�i;��&;7�.W�wc��b�C�$3C���|��	�v�(Cw��h������i�Z=�ɝ(��L�l4��T��h�]�+p�$W<z<�*$�:2�/P^~&/��
n�/Z�0<\��/��?˼1ͬ������ J�T)ɀMX���bʩaB�@�����H���hY�E�J	�
�EW�x�FJV��m�~8��h�=�1�J=*=u��R��p��\.N���._��[���IPS9G�{��O��h��q}�0P����V;U������{�5���� 8��6�� EA��X(J��� ҋt$��Rt����P�I*����W�% - ��I��s������ˋd��S�羟��vg����+Y�����F=��!^t�ߖ3��A��S3~�FFد65~,r�)�O��O	1Đ��q%+�U~���G��ǻ&i)��²,�+rX\�{���oTX�\~U~g�M�3�lM���r�At�{�7{��wDȄA���G��GђS~�S���]���mq;�]H9�A�8v	f9^I�1�WO^RZ�<�bs��\���\��?e���� ��:b�S�YB���wO�k�◉=�)0���n�K�Q��S��̉�J"��YI��C-S��6�Q��D��z'���Y�������,6*EN@m�g"����N�os�N1�]w��yY��օ��ܯ{1�a`YR��d!�]�R����	�~�V�ｇd-���_uLl��+1��A�x?P���E7�kװe������g����w�k]�A^���)˻a]�����h�fo�Ж}���&����h���W��-eT�rN��0+ߟ9^#��1r���vCo�B�]���T���&����:�f���K��ߨ�����K�~2G��>�"w\�~��㕡���ܨ���G�$�t�7?��g#%r/��+-G1j�=��f1��B7��E���#�Eϴv�&_ύ���XHm;�/T�čs_s>�1 MkTt�l�-��y�lta�\��\ ��q28�1Ja^��V���l��c-��1AoB��9�9��{���I ��.��q/�ιj3��Fol�|�)�y.B���P�է��.!p��xSc�ZĘ�¯�g0k�J�����n����[�Sw��<�Tk��f�W��y;"l#'���h �W���$�J��nƐb�S;��H��DSBɯ�_��C!J+˞�W��:�E����	���*r:���<k�༦&�w�y���Ǯ+�!�O�%�m��U��k4)�D�.�1
�b��3��ϵ�'}Zλ��I��c�&?�t%M���bD�3�2�}%{2��ʰjsi��y��S��eՊ�Q-�<����Q���a�X����>�O�]���..V��� �������m�A�9߅��,f�}Km\%ѵL��'�"���z1bw��ظ�둟n�uO��d�!	�7�[���۴3��������핪�ɫ�T�=�ZQ�G�kU�a�غ�ۃ�לB�J�l������:�M�JsH������<!��5$ka�<vc}�k}iBU��U���:��Q: �O��);%�k���a^ZŲ�'ri���}g��=M:�d|���~��	�G��q%���!�N�m���e�4ks}�LVRS��jֵ�F�x%zfﰖw�p��}�Ő8�!x�8z9�C���)��H���<,�N5_���}�U���Z�{f�1_��Y=��Kм�(�Ŝ�؏���"!��~_��9�`ۃ�;���z>�K�J�v���~�UFEԅ�Y+v��Z�e�X�;����4��$�/�ߝ��1���`{���E���Ыv��~���&Ԍ�4*m�?�pBz)����
M�*$�!���0����/-H�tۛߋ3j����ƞ�Zۦ�5���ݧa������?x߆��ٿ7"Y#�t�WZ �TFX��������;\f��mB�i��ά�}eg�}1�?�L�>��P{x��n7��M�#K:5f�qB��m����xr"� &8{g�L��i�e���{�u@0宁���jGƐD���֧'T��'ϴ�J�?�=�{9LJ�jԀ�a�T�> ��g�C�L�WN�;^ñ0��J���L��ĸU&�W�K�Q�ta�
)�Z�s�C��3[�G{�9�9#R�6lZ���~��s��ٵ��c��{�T���W9C8����ɛ��z���bo�(I$c h�,��YmS .�90�d����9>g��j�k�3�N�^�N������ʩ;���٣&m�F��t�G���j�6���'���n�U�G���q���'rșLǶ��"��O���;la�j�b��F4��An��Թ��p8�poq���e`����}�Op��*q#�?�6���wP6ZOJN�Yj`��L�V��H��6�����˞8v|y٬�>'��p��ed�i����f�P��Y0�:��¸⎠�3�����ϗ=����J:�
��a��w���eh�������aʲv)e�3Y�Nt�]y'�ʩK�\�rىB�tC=�4r:O_hUY�)�xJ(pE&Pj��8�U�z'b0��V �C����p��%��~@��l�Q�]1�o|u�1�?��j{>(�@�D����e������|��ayT����/z���U����zc�L�L����F]<�;X���xt��a������"3]y"|*-��%Cr����'p0�H��MkiP��%А���"���y���\ۊ���U�/�.��|=���5��J�CS��j���q�]�q�k>m��%i�<L~^�ȼ����/��L��w�'z4��r21@�lMV�w����#s�}����:R3�D���*�ڵ��ڱm��N�1�on��~��.Rv7��)�;�[<���r��D�	�+s%ش�_�&r2"��H j��d��\���^"y���Q�8�b���F�ԟ��[�y���˾=\8R(��AvM!MU
���K#�5��K���9YiE함�tf�}�K��,�F�@���O�Y
�R���T	�4�Ijs�	�u~�)<i[k�^\���P�������n�2���a���.
Q��V�Z�Yk^gč�M����C���N���p[]y7���}N�_���������b[-��\qK}��2Q����s�]���<����yW�[�es ��i7�GM��i��@�'��(O_�CN�n���K��T�Y<�����}��]Ŷ�<�=�&�R�"w�4�,�c��wN>9���40+��S��WY�m���٧V�5?�ޢ�0��.��₞+Gc��Y���V���*s[ɥӬ����X�&�^�1�J ,<}@�Y����П��&>�u^�5�G�zo�<�]8ϩV^�4���`^�aEP7������mR�����M��������[OM74�V�eq�q�w��3PI�[���l�~k�m��p��+v��͸�ɹS����������ͬ�A���@��n/?��=O��ݣ��A����K�����Xk�F��/�I�=V9���.���p/��y���7.�)Ё��u8�3��Jf`��������_����C$��1T�3/����0�\C� j��u�}���p�	>�w(�"}��&'f-��H�`�*�\�_�|�?񽁒�W�y�d��*&6��?�!��#�d��f��έ�h�Տ��\�����=�ִ��1��Y�X��C&F�U��&�>�/���x�	\z�o���U֑��u�'���O2��^�yo*�W�FP{<mz�n��͘2&Þ������������}�{y�?�{�n?�u����2���x�zU̿oV/��(�#W@������Z.���k�xPp���&ɸ�ԡ��`b`�~��Z\�f��G�9_�����ư³�R&�*��iκE�6��JY�D�\J/�-���o�)W�Ǉ�~㱳F(_�?S�8.qi�a���É/�K�=�6�x0����m=��}�|�T���(&<��N$8�/�"��{�!�7�BI�
��_m�h�N�s�0����J��ª��*$x#I��2��~�T��s������n������2�g�,�œ�I�C�b�TVK	�b���fL��A��/�s�Od"}A��A.W�9�)=l���_9@��P�8���^s��C~�sF)��ԽC���ϧKg��5��<=yɰ�����9E����[�%Uo�︜���Nt�?�v�<'�m����+J��웤!�|{ƌ+z=�\R�`�=�mʫy���}]�rȑ�����F� ����ض&��q��GXg�y���
���N�0p����t��9�X��E������'�9tx<P�}1*�7���S���]uٹ��4H�p�����]�N�Jr��Gm�D��&�J�bn|�@�c�ɾ=������Ơ3f���%�!f�E�%�i����xM ��z7�f�k������R-�
{��XP�*��dnO8Y�$B���}��?E0����f�"N���&�?���XX}�[3L���v.�k`�lND^�nL�B�V��-�:������u-Ruو�f �J,1ї�ced`�������{6�,ّ�%��P>�P�G���;�b׾���&�@#Ha���(�.L�xzۛg|"�fn3G��=���h��| ��V����%3E˹�I�$'a23��;�w���󂣖ɥri,��}�T�ln���J�[�BY׵�=�+�ϷD���y�в�5��G]Gy��X�ȱ�����w���E�vW����Զ�
??�����}@P��=��C�e���]&Et ���]��an�ݓ�Aq��:c.r"C���b��P��w�d��٢���.g�]�RV�+�
�{�黍g��6�8��7�j�D��-N�c�+��9��>q�2�:�ߝ�7A��Y�|7��s�^����˵�l�����IY�@�.� {��Kr�������`�{�+F��M�{�>��'}�+�Pàn`�f`�h�
(����77=��$���'\���*�D�����M�ۡ�u��G�H��(͌���r���LL�rHa��o�w�l�;ڦ����mj��v��^�k�	=��=&�b�IS��S��h��~�ș��J�?���mH�Wu�U��~���gp3h/�����a?6�Fk牳����{Z鈳i0 �����H�9����-�n�u���7��`���R4�ٍvQ4ٻԲ�Nw<!T�_o�P9Հk;���l0���۵<>�71�R��P�� [��BD���ͳ[-�u��7�)���Ώ6	�	�S�2�W��2��o~Uk�ho=V��?Fd�0ݥ�;_���� l�Wa�vzX!��\�����"�A��n�̤�:�-�s`��/'��'��\N��'pJX(����w�t�;�'X���M�,���*.�1=iUn~n�Z��?)X}a�|s+��i|}�1[,Ho	�
����-������"QR��Ak�W��a�s�{1�e+�)�p�g�mC�[C}Axt��$8K��V2p�Y�������a6���0��}�9�V��t)?#rl��ն�V����Qe�T� ��G� �_9͘�M��g�Wٶ$ήR��Е�LJ�Z&�l��	\���SW%���= p���~8߆�aaPس��4N̴��g�@���h$ȡ'w��8Ə.<;jwT�BK��|a[��H	׌dK��J|�c�ů�Ծ��+i��u����I��Z�e`H \_x�4|�k^���.>b�S��-����|��W�Ƒ��0���LÝ,�J��5C���u�\n��s�T����=��h4��Z�Y���Ч��}<쳪�ֶ7W0#����?�ڟz�b&�,���&�ڗ/_�
��<P:5�%��i�O��?�(��lK��ox
�/��t)S��@�U4mj���ާ�P`�8�Z����g���ÿ������+�^�Y�\ؘ7��Qf��"c��=���O����v���]a����N�~]���n�l^�Bk��Pdd
�#���qU�99��M�#.��̯�|�z��+�}���R���D��&^�Ŗ�9LU���L��X��5u��|� �����H�AW��"�ԩS�)Ĺ9�USl����_�i�P�iFGG'U� (k����gt�RR�J�EQ�mmmZ�V�\`�Z�lyg`�l����7��yF~��d������ΘĮ�������b]jj`����v�l�_o��]YU�gddt��_/>t\�����']`��Q���M�=�L��oD4_���p'W�} �W����m1^E�B?�����_�F6��c/�2�/KKg�U�<�[\��6��Hn�@��s�\r~})�w)ʯ�L�]���������ݵ��x�l��
�ui��)��K�o��T��^xD�M%���r��602/u���*@�� �[ifv>>>Q���L6}�c���}�h�N��R4>榩8sKG~5�9\ Bq�,�2���шZޚ+�!��f�5p��G�W��^��Z��e����]�=Z���oB�=����Q�S,�F�7-����G�.p����Iex�I�;,���@{"�NM�	�Ƈ�L�f������d�$vga�XwZ���i5����gCCC�ee�sz-��1f$&%��/�9�h:���(9ݏ���!ʤۮ �0��kdA���������T��,&RN���lf�+%��Б�2�����mu�[+P���b�_�>�e�f�{m�c�pb�J���Jt���[��/A��T�­+�=v�T2��o�`�\Y7�� �v��@�Sݏ�����,�[s��9}�a܎��>%��q��C-�kR���yӶ��X��J�Dm �<�	�e�����[Ri�ߣ�KyF5y~����E"�g�R%y�'�o�A��Y`���� �0���۲���������<+�Sݪ�uK��I(�KKA���l���*��ќ�2�� H��C��!'. �z}�S)����h�v6�5kWf�۳�g��� 5�
zB��7�O.҈�k��<��T�^�s����O]5#h��|���>4]'
�4	�iA���9 p���h�����q�'\��Û,����}��X�,ɡ:�,/��F��Gi��Zp��]Se"���Y�)]�ņ5���>w{��p��w$�D��ޜhn���G���`�f�f?%_���۰]1�����?�r˩?Vɛ���lW�;/��5X�A:�r�L��˨��Jk��|��ڍo�5�%�s̖2�R�n���'cM]��*�B��[�H�wzJ���͔@9,�>Q��ͨf�3�z�a��u��w%�I~W���Sc�6��~8h����� ��`�*/��t����=f ���c��M�~�}������x�����һQ�n<����[O�L�n�	�ǒ�?���vU�4g�b��K�)�\2��ތR�$3w����=>�D=��J�D���iM�-�iv7C�%�fU�e���v��?�.���-��������҅.�hw�s�:c@uE�E��RGGF<k^W�Ǹ�`�� //�B�5�!���۪��H���P��pS��gо���Q(�83�[E$/)+F'_ߍ��7n�஌�*����w~��� ��p���)B���j��R�+��k�.% L�<�Q),eN]�uD��-�kR�Vc8`h2�?r�.��&�0�9��D!EQ����t���5��"ŏ�Y����%�������M���;��	H؜�'l�P������l%n�	g�:$�=�Sd �kg���B�Tm<r*M D�y,�Y#����>ϥ���%�0��
�ݥg�Y�������sa2j�J��U.�@�ֹ�cz�s�S������m<z�T�ұ�3��u������-�E��h�Oc
�j��X?�1�|�.�� ��$v��ڙw��(	vHT/}��,6��Ʉ"}��-ݚ�ҪP�W���lF(�x\ڋ o�{��k�$��-��5uxX�{T��o}��L)�]A��Y���;G�G��(�Ӈ�w�?4�����͆w�^:m1j��������K-�Εԍjo��F�f���t@���F��?gW7^�E�s��D8(�=:U��[I�}���G"��#@�ν+n�CP���μ�z~�jW����ڭ��=S�s������gE]�6��q�����T�������쮈�Zl�qqI_��;�)�J�Վ�������2C� ����݉�����	�{���M*)�*y�M�[?�)��[��E@-�7wŨ��5�:�]���%�QC�V����ms��� e
e���Q�;~|c��O�y�9o:b�A7�'9�A@�6a��S *�ox4�<�'��mʾT;v����5܉��7��פ����ռ3695�5>>.���J"�o�n��qRq#{��V�q��*u�N��Z�XDH׬�u���+	x3�ت|�L~�`������/'U�EsH%�VW�����@/��I�J;8��~�Ў0x�-b| ��:Ǯ���	@�*ǔ��H�$n�j��{Fyi�3KjQY)��ȏ?n.s�D�Me��������ڝ-�i��%Ƚ�������Q�8
�IB�72x�+ng}5��:3���cW�-V�W����ȋ�yȴ/6%� �ِ?9�<��ߨhۻ�hX����6�|Z�R�2nW������0��i%D����O��L&��s���������.�Cp���WZ�О�2��h�ll�n|+��i��E�'�Y�Y5��\T^�m�zK���*��n�B����;�&���p�G�f�
��ᨆ�S�#�f]�M=�{��O��k��4�,^TTL��ai��*cr�ߕO�X�eɊ[�C*�n6"���l<v�a�v��c����~o�]��Լ
�zp�ޡ��~g,3C�����R=�7��
��k>Ԭ����Oi�h�F׬R��3y��_�n�Ta?�5f #��L	��Y��GCFF�
����	���F��bT�z�^�� 
�BJˡB�*紂�.�F\��UJ]�?�`��[���`��GO�
�\Qjj<��9�}e���f ��G�`�B���\}��l�\TTt<.'_0�jv�{Cv삙��a�Fnt����Z�;�i����U�B��\���VӅ�KQ	Pפb�.�a��gv���l��:���zi&�'��]��4�t��m�܁�\�
��{��;����\��sEQ(g����K��{�(!?��И}V ��0�Z;0s&�j5�������v{��+�@�{�W�䝕@�h���opD/��I�wft: ]7�kdǍ�W��-!�)�.�&�wĔ�G�ݜ� @���jݡ}Sl����ޛJ�S�6xr� 8B]u�P���������i`�ܩ_]9/��:�t(!j��9/Be�/�6g::�������5/�+b.]W�,��T�?pojLRf�Ϻ/${걺�$����=�ӡy�� ?A��e��z��W�ה��8!,d�]�A��,u�2R>yM���#��P���0HL��K�Ml��S���wܱѭ;��ԩ4x���f�-yH�r�3�n����+=m9w�x?@�JGgPP~���n蟥>w�-�+&yQ<��$����s�z�_�PfX�z2�N\�kg�1�WD��Eyq�T��!7Y��`��
��ܣ����
¯i5�<lJ�G|�UH��	�&*�n�(� j��ChK5�_�5]����VWB��Q�ą��/���o�[�A�����%ƩD!;3ڡ���E_�Wb�tn`�]��Ǐ�>�###�8;+�.Ι��������·[� �j��S�=!�U@���_�f������V+��8��j}Q;��T�cP��)י]�S�	+��,�@� 7&; *�
ei���9v�
���j꣔g�;���ęJ�H�R�\Ks�1�ąM`�Dhʽ)+� ��F&�;lƿ�|�o�
%ˎM�ߧ|���t����W��w���3�jˢ�g~F��<;�5����|�� :,^�7�~\���F�5��p�&���.{���f�3�a�-Qqs+
�H�d��5�j��
�>��`c��m�+o_�0	ʨ��ni�K/S�?sE ����:7UͺƳjj����y1)���V�,��Y��٨�RRR{�ϨE�{PAz�?�<��P���D�X�#�(��q��;QMI���v�� �X�ڂv��� -��j��w�-�җ?���K����rF�sY���_i��n�\�ڷ���u7�w?��I��[�~���t��1���݅�v�V;��P�?�_�ԹT����M&�(�E,�"y��w��E��U6�� 4�ȱk�{0k8Q����V#�����WεE�5Z��W3R��ڛ��_�^�
7n:u�/ �R>2"lj|k��쨤h���b� ؜QSb?�v5 ��>��;&����x�~A;ِ	�S�~4�}�C���@�sG;��э�PcGǝ���35�]-����ӻg��я��a�;��{����ƚ7�<� �#��m��fo��tDTTvEE�PHbé�����h�C�e��掑���;���2��ўZX�2�7����ٳ@�NL�q�6��rU5���c]x�~�2�'���l�b��镋ўk9�M<2-5�bMr��e���Jƛ�>������˒���y�J����9O�Y��ȞW`��!��Q����Z��_��;�ʁ4/�S5L����{�1mȷu�8��]�"�S


/���%����>��m?G��5�}o��Js�H�SƮ���:���?��ey��̦�.0~���I\�����ɩ�����78b����hk+����F"��*��cV���HRRa���?���%�� ���t��h���$�:��H�������Z$9wWJ/��\{�G�+j	v�d�� ���*g�غv鞿j��*�h����V�@�8Ea*ٳ�gu��?6�n�O�O�;::�f�e��w7��6b
�Y-��G���C��	��v����x��K�n��UU�vɯoN$����kG��~� A� �Ĕ1;[[�;��;�T��ʤn��'����ʺr�F�X׫:���x���tΟd�������.��~�{l��l�=��$�����ҿ]I�U���&�̉~��V�9���^������`R1uS\�����x����fff�Ǯ���L���"18y��4"��.M������%���ˁ����)f�X_�ߪ���9PZR���<?����[���YS�4
o���;;?���q�M�8�̧׋T�y$;8:�?;̫���P��h�ԥ5�F������|��w{?��������՚)9�\������Lܕ���EFR��/��z�鎂"v�H�����z{{��mm'��2.;ű�D?���TSS�a��ID�FNrh���0��_&�3�)�����9�[T��\~�~e�A�������ճ�6�<�X\�� ��������~��+++*�^�S����k����b���]����[���dx{{g����`�����/_ڧ��E��ʿ211�E���}�c������"��! m��;����&��I�Y\��ot\eP�����\Gg�+��x�G;x06�aø������Zz&_�&V�Ԩ���H�;��S�H������1���%�����]�Ȉ岴����h��c��ס�\���Y��㳓!�Ԩ1�����f�/jd��>��N pE�NqswX�O���.LMoz�|,v$�	m�A��"v ��YI�P薔�f֨��M��I�!�
���Y�m}�"'�$���������ynq���ak�Q�_���p��WLe�����hhh4�s�u�UL�NPH����O�P��ˠ6v���FS� �;������I
�K�`���x���mY�hSɃj7m��7o�\��R<��;���NO�`�LC��
����e _�D��S��h�-��Q�y�NIRA!�}��*RSS���j��aB|��3g�8��9!*?�1�C����F`��Й �9�:9P���|�PҠ���.�2�� z���O���p&�u	�o��k�������������
�-�@�ONN�Y����cgg�+b��5�u�1��\���������;��AR�	�A���ZZZ��`�F0>���5%9�Bw�a0�\�⨧בI��_������`��~� ���x�,�XzJ��";�\jw�P���!z��ӕ�(��"oaA�X�򢉟��'ii4��8=Y��f>{���&sy�%KG{����>د-�~��TQK8�2ޟ�VqE�.�m�&t�(�߳5����_U�$��` �%��Ɋ�8A�5t���S����z��������;0��a��f��pC��a��� ��l5�F�>�3/�� ��,A�D?��S�W� �����H8V��<��� ��CI�U�������YM	mO�'����ǐi������[��qq,�9�۟�Ė��e�(��k�7<����Q�,g���|�+Ն�����{����ERJJ�_d<���秅@S�r�T��1�2�&45��&4A^���i��qE|���#P"/_��*++��b___T�$7�`���6-��� ��(b�Q+�JK�, �c�F��cK���2����;r�K��F��B�_��'6_���� R����I�UU�����EA�ei�ȭ|4����Y�봋���tZr� P�M�<�&�r.l~&�"���)���&&�v�/��Y��3�
���_�x߿�1=�0!M	��������|�xh]�Ǳ�.�x�v�'qtO?mJ�-�|rH����9�RuQ��)�!�+PM=�����1���h�kl��4��uS� ��#�\\���q�c�y:�Yԡv9����B����e��`0��JO�|�Q�����+���k H��O�@�h5܄�+��Ç0�?��NHK���jS9Li��)�Oq��Y���w�q|a���p��R�{sNP�i����� �g|���:�CE�\Md�g��]���0{Q���V��)�s�da���vU���u'� �XF=?5%�����+�侥�A� ��MZ����
:k�=�i���!t���H�R

��5qo<� a|��4 &n�@$J��w�Ґ7莰ބ&����ؒ��� \�;���6�6����X���ل������ƺ���'$$X��j'�=�#k�_���*y0�cZ�ӧO�����D��uv�~q*�Y�-ѡ��$J��sss�-���;�yM�Q2�BM�FFF�>���q��b��u�-���n	xp;(�M榦�� ����~��3!���.>,�ԧNA��b��=��W�X��'< ȫ-����a�!�
�
�"���Է�xyy_��l���䢣���> � @귾�Zd_��/x�˩�j����vJJqN����mG���~b�X}��R{o��ϸHuk㧮���r��B&�i�����(�4:#���=ҺR������~'����3l��b1H l`�b��c�^��s�:Н¾���ﻎ��TF��^��Q����m͚r@�@����<��h�eē����.����*�~�aB@A��EM�4����p��*9ɀ���D�Sp�83�A�r�Y:v�lo\�s.�ڲ��7.���Z�V��IP�='�6!*�ӕ���M��*s@8�W%@��Y������\d)�5d=��jVu���ŋK+�����\�j�(B��^__�z�uĊ��|��['}B�����w:`���
��Q �\��L a_�-�*��]bR�ޤ�� ݀Y���QO04^�V�z����XZ�������K������P��O#�?��%4%�~�ɼ� \㯱NɣBw
��~��v����X���m����F��m���;�Φq����� ��K�ݤ���oV
.�z�-%�߯^�� �.J�ռ߮OVi�n5��j\��J�,���&�ӪDB���}�	�d�U;!~�3�x�E�#q�kk���� {�}��fT� Tt�N����g�DMZ�ݞW��ߋ��M�6�]��
�P���њ�[��6`��K�ѿEoU�QŔ�]�c(�b�iaT������{[EM��iS���^�����U0�ʗ�Z �`;�N?�����^��ɓ�j=�su� lTy�ed��靉p��ē���e���L�Nk�DW�ŷ�j&�Љ�3�)Obo���N%{�F|������I$��N�WC����-ܐ��)��^0�o���MP]�6�s�hR��4��-j �`��4���;FO�N�n�3����(�3��D���53�wjJ���۫*�AhAEɚK��-Pb���Ф��"�������!@DjHLLL\���~I*�(IK�@b �D���iy��^�]:���A�T~UUUN򷻥&;f��+D�u1����qj��/	������"ٳU�@�N�T�vV W���PB����<�;�Trg�����?�3/]���qF���o_�|9I�� Ǟ��@_6-iJ���Mk��;��L"�5��(Oh��m��\9;� �.@�hKx<�Uմ�V\��j����<t�P���\��Gy��#��}kft�+'�������
D-+v���uc�9(�s�,O߇���2����f=G���.0&
��� �����_gń�%�=��D�^�<CήM��t�h)Խ\����G��<H<��������"k0�#��T�޼݁�����x`�̼��E��#=Ӓ����k�Y�6 �@-��ń�j�T�	vw��8%ew�ƹ�dPO���N������K�Ɛ)�mN@�UH`x�����zx�^)���4G_��X1%Ya�	��ۜ��C�L�R�a.7��)�T�����P����u�D*,�|QUQQa��	um�X�?��C�n�z
���z-e����H��P����T��({�z�MW.<��}i�2@�3�-�3c�Ы �Z�"�}��y:/����#��ʊ
���t��мV����������ԫ�F�[�	>=m�R�7�����sL!z�{k`J)�T��p��X �R�����������;���`s�a�E�^�+�]䕽������L����1)g����I���k�j��Ih@'E.�ZZ�Z�+��x���1�.)]9�.���?�LRڨ�OP�HyG�+�w�~C��@ *Gh0��
d{2	�Y�HV���t�N��V�|�^A֪��K��G&����W�̀��|�v��{����44rY7�a(x߉q�~���O�)�?�T2I�����.{TH�S�x����[[�&��XGʯUg<��)b�� *şj�.*�4a?Z��/���ʙ*�������������m�
dP�����p��y>"2�!�ѱ��r�l i�~��y`HEU��6�������]�}��vJp8�������#��3� ZЦMD�&1�NY����d�~k�Q��t�v���U��k!�A��x���nB*rR��xd��
���s"��V��Տp�f�>����D�u�� ������J����67�}�U�e��)gbV�l��(�M/ٖ66g#��C� ��c���x���n���9���ꛌ�>�q��G�vvh/+I$c.����

�}�:C��0;� �n�	��?��m��SKM���y� �[W�׳ �zu&�PX��r���`N"�詩��..��zZဏ$i덅n���ɨx�(Z��x2E�s֚I^�h�&�I;#����ј�Ud/M����͍��)�E�^�F���K�GKS�r.`wKY���Q�z�h{��?ۛ�@&��줜Q�ܖ��D+¯���fg�
�}*SRZ� �"1M	<wK���~v�6�7u������џ}U���СL@_U�iv�/<���j�|Dp�-j<]�>s {(
6@e��)R(�

�*��@�����B���j�,0ߡ��H`y������)(�v\||�:|���R�� �R �6�=ڴ9�y�����'$X�]�j5�	���јN��2]��Ӫ�s*pp=���8
i��H z⛣�iK���?���hV������<8i*
���Ot��ݤ/�	�m��d�FT�7�|#�ٙ�@�`v��Y9�	Í=��oۻrѢ&O�h	\���tM]������NHS�42-9Y��ԅO��C��D"N�єf	K@ ��T��0l�����mq�ͥJ�t�A��	TolG+(���q�`��p�Q��=.	���&� ^.��vJi-��@�����u՜n�K���ъ���J���c��U��q������c���Rv���?��ݸd�M�\Ԣ��vŦ9�⊻�[d2.>��f�׮M��F�ܧ�n津���鎶��v	�s.�*(�*�oo|~Ɔ�	�5�-�U�I�z$M-�<)1 ��W)2VѴn]Yh��4��������u�pÿ�h���	����n��'�	E�)-��{i��m��<9�]�->ƭM�0�@]�򰵷?�Xw7��A�����wT^����A�L@��j�٢��y��6X���{Y�8;���2h9�����	P־>���;�w#T
�"�%遦��xW�S��x6�?�{w2�l�w4�V����H�=JBE����3��S$���S���כ�ii:r�4�*e�&bC��u�"v��U�Ϛ���]coӢ���q�ߝ�)c9p�+:\�?z�YC���z� J��e߼����|��0�v�3)�O�PO#����[Z&p��P�SR�kH��?L�h=�Z�ftr�"�������V��:m"���x<W�a���n�QO�ɹ"/��+)�
j�����PC�s�zfN����f��x&u)��<��	%vo)�������H<�
]��q���ǿq���&Q��l R)���������\��Y��K��)�A(A�}��Q�����ed����B��=��a�� �K�P�m���!j��=���#��_+C�!oB�����If�٠��6֐[UUU]W������T67��m����$��߄�E�qvIU�MO��0h��b�@͡/���:����w0	[�4����~Aql)u��\��_�
hh�H������P�9;kV�b2b�i�%I�m%K�([U1��쫮V����^8�hB�l3�E=��!0���K��A�4�����D!����c�T#���kk;D�Bm:�*g����Q�VI�<U`�ڔnӺ�d+;�aN.��Ɔi�~g���l�'�f�;U"��{�G�);3�i�������E5�.@Y�ZF�!����+>�Ua���\!�����.�t���n�:�#w�`�U[�T�5�J�
���y�0��
y����w���#n��׷�sS���(C��Wa�k
w,��x"Q0C$R������e}��a��t�U��a��0)���r3A=���p� ���������3%���ǽ��r �����
�Hs�f�����j���{V��F��&{}��1+pG�%���)j���i�f󈊛������hhf�'�î(���Kç��j͟�'����D|ᬋu���JjJp,�/Z2�#6�u|��u�>� ����3!B|�s�R���o
���:�4� �ՋG�-*�����ҩ�ɵM�P�Vx�E��=�ǖ5::��������tZGzד�_���f�ץ?\����KEc�3���>���t���~?�@]�gG�% {�ڄL(G�����ͩ�/S�>J��B�P?�(����g����>���*����H ��K5�eZH.TRCI<��?� es�6�T�h=x��O=-`���P�$;���"�ZGh& Vq>:krr�3����4�5%�`��漦�r����E����r%�gX_��Bo>�	�[����utosD ��=r�E�����8��l���O05M�UK�!���� )IH������@\}�Dгo���W�Sk�5DP��̅�&[�8�X������f?�< �x�~�ኴt��t� ��/g����:�䰣�s�O�$��h���BB�fP��� a��s���>�7����9��Ik�J���A�9��Ki0:gڞ� ��)�C�����u�c���/����`�w,ꯆ�އ��a���8|�.C��\{�ਛR|#�Ro�fNP�MZ�?��FYk\�:����p,�=�ʹx����|ؘ��qK�Ԉr�bŮ�(���'���u�o]b_����g�� �8�%�/r0Q+�p���i�����غY�?��\�L���a��������Y�{���o�kE�����.؈��rZ�!#�DV^^��0�$a�7�[���F�d�$ K�;$N:B�R�Vοn���PK   ��X�� �f  y�  /   images/96fabd4d-0b16-452b-94e2-688cfcbce531.png�	TSW�6~q�i�2*VA �Z*((�'A�0I�PQڊ"��"2�A@D �A���9�s����������f-���s��g�g?���^��ݕ˄�A����F�<�-Y�X�����_>~K��/u��A�����������t;�d��y�����)k�h�>s������mĀ�0m�j�;��k�w27���$[&f���tt��,�ｦ���ݒ�_n�1�`�=��k-]|�!so�O�~oy����B?I��l���K=�w4��؉#�[^����c�}}҂#n%�@�'�M}S�L�d;vg�|\������zƺ�WOڪ��g����VW	@*<�6++KK.��6��{��4紧���;�쇿V=漘5��L������9/U�c��r��;]�[�Ťk)�zj�]i�19I��DU �ƻ�{
!�w(;\Q4�_v��ͪ6��![�V���1���|�;����0�j�t߮9=X0�B.���L�0�C
�17��p�d��ۉ�� �n�=]>�����A�oVtɻ����1�Nj���v�.&F�3T�gČ�iL��S\\|����7=5��SK�����,�2���؟=���/ʖ��k�޻c�ׯX�p�@|TozƬ�N�Q�TcIx��z��j��xd5���:ﭛ�_��cz����5��V���D�Va	-$���E!����Z�����n�\6�^{�-��0~��ߺ*y�MJ��_����s�r���0�Y&Q�wNउLL��V8���@�%]�A�?���z"᫇�\|G�*�ς]��q�����"�"&"/��M>&n{T�=���j;��{#�-���~~~�ѕ��Fd�UD_��a7�rQ�2�ۇ��.M�H��-��y29�H�Wwg!�
��YW� �ѕ�=�QV$_?�l�m��7s���H/ds{W�z���]��Z�w H'z�S%\���4����_$����Lz켣���y����a����vD��WU���u���#0�O�qb�П9���!�������@!����^�}�{�1�sN<rĂbH���Y\n_��e}�NM�*l�1׀w95�����k�;ga�<T#�B_��zu��X���|MPb�[{��O�%ot������$�u�B������)ڛ:�F.P�9����3�4���s���,�D��Y�!I����I���0\��4�����2ښF0�K=83�jLӐ�OV{�;T&���{6��mr���n�9��2�fq'.�ZҜ=�l䣪��5��9/���ԙ�6���y*�w��,+%UF�lr�M2�]y��]4Y�)ˬ�ޅJά�)N9]��� SD�,���.����^��<7��]����))t7����|���e���\I⤌�p�+�4�m�!cE�Tc�ۧ��O�����`���4��BO\9
����NHk��<.Cȝ�#i*�y�YMMMK�,9H�l~}.]�c�����86VY�Q�榆�,���\�Ǉ:$bBU�Y��A�C*�dz�gHp�x��)q�8�;[� 󰱝��l�W����\l�G�.��+wI�l}��v�;��a
�Ӎ�Y�wVA�x�˾�h��&���@{@����ւ񕒜9KF
�-�:�U��]�V�ç�2�ko�sn��z�ah��d)����
��mN��e'*�[�rFXOX6�[�D�ħ�!L�iG����I�P�qT�G�}}���{o0�N��s�x"����Y�f���]�<�RdX��~��cz�Q�t9�H-tRv�H�N��=cn�a�f��fk���[��?��B�eΉ N�]{��&D������!]��Z�=q��o��e�~�8'Os�{'������r2�p;�CD�zݽ'i������܁�---�=���>�|� �"��5�͎�7B�=[��_�K��΋7�d������f=N��s�����0-]K�S\sXˁP\uz�����UЉ���4Y���xM=�yp�A�s	-b��wn�ϻ^n�34W�pc��Y2rEA�.��`�{C^���;UaG6hsl��)h�(�Є��G7U���d]266樫m��ކ������=6z������-�Xw�a�z�Rt7� �$�](�B���-��s�G8��YhU�� p��r��v!(e21���R0��~��z��F���VnYM����љ9�tM6{�9��iͿ��*�&#A�o�g}�Ɲ�q#6VL�┘ds_��$J`����y:o `��/wti1c��?r��m'^$m #����K Q;����ֱ{��1;J�uC0�0�{��v��h'a��a̧QJSp��W���=���{ ������q��"-�l6ȗ�2  H��f9V���
�K�ȋ@�h�
 �d�W.��5r3�{k�Ó�p'u_�"\��F�V��F�nz���CF�����}zvNMu��x4��<�5b����Ҩ�,ض,���R��˗/�2^��o�a)�\�X烠,��O�\	�����*�W��KJ���a'��d����H�4�%�U�Y_��DgK�TlB�m��E���iÅ]�Hٶ�h]�� �T/^$R� �d����X��\����^9ɪu�uM9�![%� a���M0fJ�3�:a�f��A�8,d��h&���X���dե�fҔ#ybvz V)��R!;����2G��[�'0B#Y4͛s��ϺC��@��l����N�.���� A�b��(��g�H����\U�r��ٺhONl�Y����K:�
��g��ӱ��X��G�Qn�Q���Vu�ƾ��0�CzL$�%�j�M��tG:��|�2g��_�����~z����' ���p�R��X%V7D|f��fx@^�
Ev�9�jN1���v�Td紊(pO�#���sl�T��c5��B���Uy(��&�)S��&�\�$Mw�s�zn>�	ZjêkG)��=]��wX��JQǖ��������nE�?@j�����}sa�
?ᘗ�i"H��	T7o��+�6����(g�׶s%[����圀����DS��Z��\���y(Nz�DO1hXaD�J8�\�����;w��������,É��6W�i�����e���|�>�@�	��6��M���WC9ɵ�o�3L�@a,,͠D}*I}��4c�r7Ǖ��cNZAn�Ct�ׯ��}��u��9i��
�R�B���qW����Y|��i�κ"��ۦ �]p�o��	HJ�;=ҳ��8��1�*Q�t������p��q�^9ȕ�6]����Ɯֺ�'�1tqV���"(}��H��l�0��h�0�5.�RO�_#�#��gPrgpH�f�z��`��زT�c�T��$1.��Y�( �(�t+AzvI���)?�hD|I��Q( �
++��9G��G�g[F+~����&�К��f��1���g0���G�D�t�jDG�����E0��p�S�}�]��-oQ��=BPbӥ$]�n����E�x�E�.�R?�Y�CN��k��l	
X�É" �XM6�����q&;�Z�`�������D�~w	4��<q���J�����uϩ2!���E�5��(�8vu_�q�qL��5���V-; �+
��cb��03�E��w@ˇ���1�̠�&5og�;8��9��=�N�Q��(�q������H��9 �)��|����ŵ�#r��Ǉ�z���s;�EͿ��-�PN[���Q�۶�:xF9Ҁ�
��D�x<ݲlf�9�W ��xމ��=)�<ǀU�_p"��0T8foZ����Ć8�' �U����3�ј]s" /|ŵ���6��i��F�Y�h�֊���n7a9������l����52�X����zw�0�T� ��ӳ���K`���/9����
�N����
/ւ]q~�4�ڠ���I��R�zU�R�%>�`K�e��@%UI����_������FI#��o[�z#9oҽ��w4h5�o,$�K��úW3=^0��b��'��պ9��՛���'��A��[8�����֒P���\��
q:*��WO�����5�Hl+К���<u��l@vyV��B�(��A)�ưi6���WC�����6)^�� <�]�T��:�E�y�K��DϬ�ǽ��5��;��_�ѳ��)�N�Ɗ�`�p�Ig�(y�n ����|+v�S��J U��)�q���g�H��} `��\n��;�C�<�����Xxt���,1��;eJ,��-����ӢI���^�%ڍ�j�oŵ0�mn�$�ܩ��(����wS��QʨfĘ%uf�t�a�ujR2�H�tz�W9*3XSQZ9�7A��W�1!�?#����Z=� T��'_���vd6��`����Y1��y'��;�'C����r�[΂̉FrD�:�(дTm�ZUcBgᓽtV��%�Ŗ���m�����55����mQ2�����sYuM���~B+�u?���=��}"xl�7i�#������I<=��.)�{�z'�[Us@��a�q�Ғ��Y[Q����I3Rr��D�O�ƺ�61�LZ�<|E�Z�C���2������<F�`���F��֚��N5خ&�^�w�	U���:��٠�Żkw�ZE�\�ʐ��w�����)}�	�j)��Vs�ۊ��X�ЗFRfӱ�3-���{�zb���Zw��=���͠���(:�w��v��qqX�M��|���-;������K��֖K��I��YV� Zi�q����c�|0q�l������Uº����4@�5D8�i�����6纜�B����pŮ�D�שr����錩�<�B�Qf1t���Hm�޴j�e� XUL�b�'\X}��O�
L����i��olA��(�2�~$Bc)�-�9#P�����{3��r�t��mS�#������Ps���D�΂��h6���ޓ��y��Zzv/�(��^Lb�^����0؝F�Q5�3�r�ӏY�)��S_���ꝰ�m�sCcb>`:^�Lc�b�7:ekK���=Un#/�
�zk<\Yv(F����X!�{J�����zW ��t�s����\ˎPF�/�&�(�&Oh�w��a�<��6��B�1/�'��ş	�~�rl]���0�����oA/i8��lz�E%na^T���dd
Ut^q(���M�����-�̸Q:bA	z�[C���;D��89�0�zq�!�4g��gf|uw�4�4$��.�I 4�?;[�Y��[8���9S�'�BHjH����b�pؚ�����T��1.�`5f���KI�YWԹ}�2{�~b#A�h����2�\<� �20�VۖA"v�?7�ۃ4�"��������iP�p�"@�a$;�����}�*n��� ���d��-��'���|�漾����u��ɬVKJ*�I"ܾ�Jr= �v!n�r�!�Zܸ�Q���D��3+'KnII�����(Зc'��1�"����e�
�o��0�p������d�.�)� m͟��H��#�K�9�%��zO�nS���Ld=2�1�?���<k� \�������y�����%����p��� �U��[%��g�V,�¢��m�Ŏ�Vg�E�:f�W�<ȭ,"Qs����ÑFk�څRh����9h\�*3����������p��t��|�ۛNZ�.S~;+��p���bkc*��|F!�=*O�M��nM_�B�����󲹎���[W���tC�t5@���d ��P0������
*<�L�;U��M5���q`}�/C�p[�ji��kd؛yy�C���`��$�S�[25����	��c�Q>�h���\��	�t�	j�{�Y�5]�<�y����5����� l.P���,�䠔�f������+�\8-�p�-�e?A�b��d�"�(ǫ��{u��#�J6]���pݵ�}Z�� չ.��8<�b[�,�&�K�`G�+i�ۍU۱��&�'�-lϗr8iP>�A���P軜"��Cl�-�ध))��+�A�͢�;����,��tfm!��Ť.@ڲA���y��w	p?|&��PG�&���ښ��)5�Pɴ0��&��r��}λ e6)5f ѪYط�� �0Z����p{}��v��!���[гVШ�y!�;hY���lȲ1���y���������"e~����Bз�M��:K��������էxJ�3�Y��G�WB�@��P�IF��L83�cq
�֜�.*&����0�lH��Y/l� m!hi~mry�nZ�����iƞ�2s�{�[8#]����&��2{C��y
j���h9
�I��!�f�6�O��	�=��(T��^7Y�X��i�sQ		�:��AW�ú��d��t�v�%姶9�B��ŗ�}����4�~��s�) �K�,B�_�U�?������qnv�m`��ڠ⎱c:�+�u�&���&^k�MP�z S1�w��jȇT'�A��m���|vw�jD7�@O'n��o�VE&�8Fy�+k>{�84�Z��~����������?9�l���;��^�����џ�X��	?�M�!Yǿi�㭗�s���2���Xq�R���Z�^u� �hB�}z~)��14~��F(b3�\�e�M��W�p~z-`|�&��َ%�X8W�a���9�'@�?m��9���Ț��{H�A �-���7�PkVw+ڤ�O���oHӒe=��v�%�5|F�CŬ�ڒ���-Z�l���=�A,���ه`��S�X��<�ۛm:���G��}�ټ��=]8� ��N�e`IU�l.��c�hp�{����e�d�Ѽ�A)p��[rΕ_X��W!�����W���V�
o�ɖW'r�n�r22�Z_�o����<ӣ�ـ㇭�(ہ�ey��.�>aN�J����3S36t������cT�8�d��j����$P/1�P�Sߩ�4-v�'sȮ�CB�PMj?(�0'�����*e�R�a�l�O��=�l=���I���
FYb�)K�sO��t��؜�/?���d��G�il��ϒ���䲟Ӓ9�2u����,�E��s���6\ÏR�9���}S�{/��w	(���cЎbG,��/猋��s9�+9��W�c|�{�B�D�N)��>@���:9�T���s���J�ka= G�P,(�8�����^��~�I��f��ps{��w�����RR���0&y77�n��亨D�iE��7�C�i���&��@u �:%I�� 2>ݸ-=-w>���I�0ψ$�^����LX��x�3��M��(I���@+�J�>����Է
�Y�}��wKj�9���z�Ϧ��x�շ�2�Bt���
}�����ث+
j6�6��!�#�c7��ى�YΏ=��څM��*�s�������[R��쎇�:�Ŏ8'���|O�w��ʋ?���z�H�<9�:r�1*��ͫ�Z���K��&�{���~���bK���Ǣ���o���t��}��I���~���r1��M��BC� ]����z�s���4�� ��z蜝��J�L�}H�5I\p�N]e�U4CZ�f1��cvGv�4��c��B]�i���p�->o.��fWT7Թ]�vmfˏp��.�����I��qHPCj����HS�'�zqv�.ǷAj�}aF���J��DχzAW���n��j��9���d/����;3�j�H����<QA@��m^�΍�M�H3`�}��I��̦��ר@�J���ũ'XW��Y{��f�|`�=ˠ��t���-�2�r�`�0���F0ڌTz�Qs&�9����T*���A�i���=�$��P�ej�������|dl��qkAzzd�>�tU�4(Mk�48I�4o�Y��y/�GWg�]�Vp�I���P�c��%_��Ž���&���$��N:�ň��T�f��x0.�b�َ�m�Bo?||�l��Lv�fsj���q&j�2gaFeNP.�3-=E�PSS[Lu��el�x�U�G��}������e �؃�<w�r{g�-�op�q�����p��н�|R�*k��܉�Re}�n~�.](�b���"�7��΋���?��.�A�n�ºu��Gkf��0�ys$�ʻqL�UEa:��^_,(b���`D�ǰ�@^�M��\6�V4�xyqJ�!��Wp�R9i#����%��Ka���?�q�{��� ��魷�4�[����LQr5rb!�gÀ�n��n7���RDӅ=�,*㤪Ho3�7wgL�|.�(�0���!7U��`@|�e/[@'bz3/��2�Ҧ��ϑ��Nn��������j�R�c��p��>q��#c�hE�=��_�@�Ϊ�Jbe�?YPn�R���K��Ka�$W���­�I@90=pYP�+z���ƹ$Q�����J̪�Y�Kf��Fֲ^�dj[J�fC�K�+-�����:r�=P�r����Ĭ�E�=A[�eZ�P����]��4�pJWH���4LS9�49���5)5W>E#~W�A�M��ܡN�׻7UMM&�>�P-��X�0�q*��~��k�'��)��^Ajj~�D����TMu)Y04��4�`�aq����Lſ�D���R*���rnQ��	z&P,�=�������{�#���H�$b�@���&gS������1S-gf�Dʞ�	���]����	�������=�d���\�?�n�����������������������������}�.&F�?i��]��@��=�ֽ�Q���u�e�˙а�K�S�={����L�ym<�8�+!��B�qO:�;)����C�#�7j4G�$�I}f�M�K���`eb�Z,�G����#G2���F�&��뭣�X���!q�挽�~(��F˭�	�k�*�����Oss����N��9�6�����V�xa痼�����h%��Ω�FM�P���ƐK�ǐ����hh��Y�Sk��Sr{�ݛ{wwe~�c܏�n��d|P�b�Ӓv��2g�<��}�NIL���=PlK:�tAe�@��"
�>�u��3,�,�9)�QnsN)"rʧ������gML���ه�:��z��?��r�������q�/�i΁�w������[��ឍ�>���q��7�{�_ޘǬϊnR	PX��P�;��ҕ�5��+*�eC�N��]��Uי�{Ϸ�^�s6�]��M��-R&�:�7��5%;�F��q�2�e����%>����}��,�#Ci�}���K�����K��@C�i-�)�c�=�T�;��DȐ�9�aR���G�a��C!�M�N��f]�+�\�Dy�vf�BH��$�B���ֶ?�2�);]Nz�KIj��A�N�ZagF�r�B�i>4��?zo��Ջɋ��v'�F������
�Yu�+�ϔ۴�T�MLu��qvf���ʨؤ���x�>�Ŭ��
���{&�Ns�������� yG�@�|\\�����sg	��mf�ŏ��Ë����@Hq�G(��άoqs�e���h2G1����K��GK�Zf:�h�9��b�r_�ϫ����l�a1��!�8�}gggBL��p]�&��o����dd��O��o!�����	����@>6��M9�l+�R�r���t�����5�gI�Jc��������[S�\���X�i��
�M���*؜����
ͬ����
��DV�2��Z���di�(Qa��|��+�_�ϑ���b����:���w�����
c]����'��`��8-D+1���D�l�Gu���t������Kjy�ZӃ�}G{jz�C��`{Q`��%��x�.o�l� DX�r���	�%kwӠ����?���͇�z(��N�2�A���j��~�]�r�o��SU(/�'̤�ncA��:�O�Մ��?�*[_����G�we������o�v�X'�
�p�W�d��[\ބ
�( m���:��g�c
y�Ajq���%��M<��'�D����@PzJsV�:�^M5َ󯣃U	"ZZ��*h#��"���V����+)Dg�!��h3�	|˸����0V�2����*~����KJ
���R�k�7݅w/&��W���!������);!����
�z�_�m6�H�Z_+��n���λ>"c�|�.T��~.�kV�
���Sn�ŤƗ1�m+�Gsn/_d-7�R~9�O���m6����� B[�W]��-P�a�"�ٯ�η�a9y�u��-��6�\
Av���< ڴ�)WZ[F�y��4�T�o��b�_���	��#���ԻF��I���_�M�v3�k+ hծ�ry�ҽ[ѓ������n"Q5����ȷ���`�5�Q5���*��� [1�?j߻�Y��'���%���m!�91)	9����k+�P�"\�[!�{Q�������󡽚��MX�5��4��y2�G�������شC4E%��'�W��dM��J�Mc����׈ VΡP�W� �y�J�G�,fm���W��M����u������9���+���NP~�
A�G�w�$B$���)�������\�OW,�p~�8_⓯��_������_S�(T*�� (�%o!W� #.�R���s���t� �����s�x_����A�'`!���L�U0f]��`���J����H+㚗��w���S��.�<m��$�L@��J�t���L�"3��Oa����(*�Ȋ�����&����Z~��p	Xi��1 ��o�C�_q&���tij"h*[P}��FezO����X��r�K�׾_|�ja]���ѻq�YOц���.�:�A2N%�hVs��}�]����C��T:�˯*��O�7\�3E �(�ׯ����c�������t@�D<�^J'�9�Ci �<���V�G���ݹ7��U��X�������j@y���`<�!\��^� �C��'�'L���,�OM޺f�B~Ś��?~h�s�\{��|1��,�������pqۨ�H��0N�/@�t��H
=v��������d�"���[�������߉�K�|ʎ�?��Ż�F �EF��o��q��0���x�����5H�2�}n��Qa{/��R2�Ex3�>�+76�{��͡FC��ٜ�����2�U�?�/�����Ĭ��aS	��mF�N@�vgtEL���7��B��������� �]����߽�;����Y_��qtnػ���@�j6,�&�cU�ߋ�'^�k7�s�u_OO?�s�����Z�C!Z�Q(/n?���ۡF�w�&�nE͗M��F �J�Hg�{��G�@{� �ٺ�3��2�c�V����$�T���~c��@���>�6%%�0^W�r��k����ZS��8�oK"��NI0�`�ay�g��Ъ��o�}�n�\�6~Ϸ�M�!����Um΋i�3�+K�c���ʓ���������T��K
�廇\Y�;�����3��-��X��쒁��ݠ��������� K��ļF��l�H[�vgj���;-�(�Z��˩��wF��b�O��t�(\�14~9�z0񋔆�`���hW#�LQD�y�����N��
���o��maN�,5������6�@Z��ֶ������F>r�?;v�I�՚��|�#̛�M��J�
yvƆ� Z����L�]�l��i� �{��z�v�����V�N�U`@j�������s�d���J`���L�[Q�\��Z����3�B���嵴�g_\Ӻ��������hÞ�وЪ�H��+Y�<ˣ����$A��{�ױ��ة4l ���Q~��I0)z��#˿V��n!�����d̚���4�G�k�>��Ą�ؼCQ<8ǅ�����k��	�P�v�p���FLL<mwww���
�L!VXQF��-���1���L�]�r�H��5�3-h����0�.�5Qr��~D��Ԯ���դ��2<~8'9�����d���qu�� f�y��WA"fH*����w�&��.����s��!���ҒJh���ҝ/Ȼ���nnktuu�g^�#��_/**:ii�y�E$�Uxb�S�V�M����
�� edd0��>uq^���`�S���0�1!1������G�L�ə=[5��笉�/�_�bl+�<�=ݥa��h�F쐕��W9�p`pql��
㔞]݅T��6A���cD�HL�e��f@Qnb/�콙���i�)�!�(+RE%����^���%��4Co��j�cZ�OƓ �͒ͯY6W5�V�vy�G�?�Lu"�֎�y*��-4ճ�32���W����H����Ļ��&�����Ӵ4���w�?o�`PA��;:ć9(�#{wz?f��h~���
#�j�/��a������mll��!�~��.c��[RɕA�Lv��v_]���jޔ�������y�ӓ�!#<<���f�u�N��ț&Ԛ�e�g�P����X�)��4�_�!a�F���>�J`NS]���79*'Zd�	����Y���b4Pv>����������Π��(88�د]Y����v�l���.��LF~�g�_�g"��]L\�Um�	��������L��7=�Z[]]���zݲl/ě"I�I:4����W�^��[=��X���'E�b��3�+ ��V�T�j�_���N?)���c}���p��H)"��x�ԩ��1�'���J����Qߏ�۠P��
��l��ɧ����Jt�2rժU�Zr%V��°�����'m e�>�s���:�C�{��wQ���]N��	i��W�H�x_JE{J�f v����������>��Y�)fć<a��(�3�n� i��6�b0���-*_Z�����L��kaD��lR6DP?<B��mI��5C���xQ#=���. RGc07I#���*��̞���-�Q���>��(
u�А���^&&5����3^���Ky4@����D���c��@���=k�/_�4=��[v�����Q���Rw�Naˁ�,Đ�^wf����&S�<�.^L&���i�ɼ�� 0�$Z_e��]���]tfp��;�HT���5�t�>�[���Ei��#��.���(/+��~� �w>�Ԗ��Hۜ9�@R�]:^� {�d	X��4�1И�B�5��I'�������X{G��\��Gܲ��+
[e)})J�|~t�p�ATDdd�|�,m1L̕�N�j����d�j9,C
3��[�̙b�SB����]/^�8mo��^��99]�(�F92�%8 ��T���]�� ����ʾ��m�+<��`�U���3S�/F7 ���?`hU ��ddWWW(S��C�2�6e���dV���T ���Yb(TQ�=�Au7����툧�e�ff��U�ώD7�{�	����j�5xO����pU���(��熝�K h�v>�lc3u��G��`2ГYY�1�K�SBR�P���xt_Qs����P���� 1�Ԏi�=B+����x'���
��#�1�]u9��b�mB�s�$m���@m��'OΧ5Tv����NH茏�$�s��Q<}�Jk Fh����L�u�2��1\MD?'���m>$�2P��<sr'yy��϶Q��4�@S` �*�"�s���'��3�)�M���Qvt���r3��K�ݵ~�I���m�,��cH���㴭����{�D"�B5�l��)2qqq���7 ��D�@|R�V�]�l>;ҥ��W�*4B������J�B��R�v1I �j�ʌ0����H��%˭ꦬ&GE�$�#����c0+�<��%+}�w}��{|e���T#�Eu���������⎺����I	X�?
�	�����5]�'��0��y889��O�i*( ��Ў�	�5�kIꝌ�+C:�Lʹ�z�e�ڟ��@@� �XP\��)�A���T���Mh��l�� e P<����#0�?m)�(,Wn��0s"��̍<���l9�BT���p;��A�&SR�y�f2����������u���!��S�"�\"Q<3��,���A'��:б�o����M�(7ZМ�6�цdp�L@��Nar�9���BR�I$��xG��1��,��i�^7 vy@:R8h�7s �:Wr����cE��y�e�>q�y��S.��5�;/+ �OĹ���j���a�n;�]�����qfgh�v�� @�%d�Aѹ	���$��E�]<I�����'oe&2�^�d�=I��T��x�g���Hs�pQ�该21��xV�i6f�E�����ˍD��"a=���Ǡ-�*uo��BG�,1�_PP���~󚠄N���!"B�Fjr��N�|���Pt0p7�u+�$E^Aa5`)�]P;�aeb�RS���u^�}Ro&�i���EBi����s�+8X��+B�l9��:�:�'OI$����J%8SZ&	E5۹�?ाLBL(�e��i8��#c� 0|�4�[��� ��
����n[�-�ߣ�0�@��Q���R�*�ng2�i ��=�|�_ ����1A_Q�O�'�,-M0\�������ݻA�Y����M��D����쎕���&��清���/��F+���L��N�N�Nk�,--����G}í��O�4�=P��~�W����b����ک��z������9�&}}�����ޢ��;���;F��23�{�XR�fW�ׄf$xN�:��ȶ�ZO�	�#\��5�5�Zx�$�F��Z�Ύ&E�\8��/�ٔD ��ڀP֍��XP�����^��B�-�>u����A:��ҁe��I����EnG�b7���HH����h���G���roNLL|���r�`������_��i�SQ��K��u�{�,�<�LN��&��&��=�O�@��>^��3~Ƞ����quD�z���ji���O�y~�hr���;��&Xao�篵��C:*�u�}��$a��<���/_���y!�6QX����ud�&m��REEE���M����?7M }w0O8��,���mx�>d��a��W��;
��O����jۣ�XC������8��sF�u���Z\'��E�4қm�9IF�Տ�@3I�o�G�����#-3^y�GQew�p,?�$)�\�?�R��f.��F��J�:L� �_d�7\�ag��|��u�C��l �<�a��k���ƺ������5�6�ު�ݱ'J�.���U���?�AxC� t��m?mrǋ�u����(˓�^gl5UIA�mf���	�?b�)��`g&{��t,����1*�
ᎎ�! 2��I�Ɩ��&�l�̤�V�v�!b��l1�+K�2�<����6�0ةP�8��l>6��>4$/.!��h���r���9�"ch��a>L�`X�񾊢t�gq���4�l�ι��Nͅ�	�YK��h�V,oHC�pe1�v�C�ձ�m��A�w�����o�\��ݛ%<Q���5Ђ��/��-E�K�x����CԧMJ� ݵ�ӫ5w�W��,:��>o]xw_��"���މY�V�s�BS6�$oe�w����{=�'�n^z���\`��T��O������K\a>$���K����S�6�*�yVI�w�����z;�	��[���I��_�w�o��_�^���;+.��m��χ��R{��@�%��!���=<��7�@�%��&�D�'�Hֶ�6�F�M^��u����:��c��&�/?�ٶ�f�N��p(؆����<�p��M?��]]j��}Pr��dYQ�|]�L��3|9r9��>p�0�A��7X�]���o�y���V�q�+%��ٽPr,��!m��v-�;�+[y��~��}}�K�1���hyz��H�8^[#dd������@�ٻS��9�`��;��Xx��K�hn#��_�� �;��ut����g@���ŗ/�o����n���o������?yA�)�
`%<�j5kk^�١9㣹�-�ʧ�o�����@�������y��e:_�(S���H�O6>�9���Q�{�o
�l|Qt�n`�����0����7��pk��n߫5
��}�a���l J�������,d�8H�����AQ�V6Bz�������p�͍�]B
��y�������̳�� �̹G��_��S���>�_� �D�η����T����I\�u��
�S<^9���|�`:ߏ���D<�}{��.��W�����t���n�Z��l����*`xy���!6�_�:����.GȼxiΦX�6P�&D��� �� �V>쇜ݬ�y���0ʻ�kUa�p� �R��v�ڐ׺�K���E�������${������zo��m�|N^����9�	�9%�����d����ޡ8b�f(�[��{>�<���90������r��i%������_�q"��}1Du���'�]yf�[�K ��;ͣ���8�2�]f����jcF�c>���������m���"����W�8�Ւy�ڈ8�=�5� ��Ȃ�)J���_L��y�N�l�S�۵�l�w��+��ϠA��Cbu�^&@�':���qq>�G��?jȤ�W,){]6�4��Y� *��V��&N����J�q��:=��?���'�x[DӏM�z��������Sޔ�{H]}j��"��_�DxG�O��7W}���I�Mkxt��Z���ew7�a��eu�M�dRݟ[k���H�o��}V>e֡��#��>6�>���ҩ�oӾ�<=�b�J$�M�K�\�Z���?�-z�]a��I�(�y37��{ץT�d�����W�/y3�
s%N�4b����t��<t�|�v]
�����F���TxA*������'X�=x�ܛ,�k�ª�yi+��$����a�û@1_AVm�~ H`�O��N�C]����G@���+@��%ށ�>AX���ޯ��OQ 9�Lɲr0�ｚM�_j\>S�k��9�|�h�I�d�����C.Z��2����]�{���E;��}�e\��L��x�!�BGy�h��s�T�'/7C*�G��Nyx��ٞ5 !�/��|Z�Ma�B����ޏ|�anT�2k��	`��_kƹOk6���n��G�V�/��7��b�~Ee�E����BC�WD�����^�ֲ�����6��{���5�������ξ��(��ln��	�D�1�)t�Kl;i�� �n���#`�Y�dz��?g�����
�
c�ྔ�/�0��/;�?�$��l	۟������ѱ��F��:�WF��6O='�k
l7��>�d h�ꗐڕ}��_l��f�����>���F�<�����u���S)�ˤ�ӝ��!��Dj
PsC醹��x��E���A�;�8�v�%�JA�d��R��
�9zy��ҳ�]���s6�������r�B�~�<�q�~����O�QV��7��9��&@���%g*����kW��]���4.��a�`N|�;�H����~��$���?�R��ħܠ��k���̗��ؿ�� �`!�,���aF.�ka@�#������O�#> f��Z�|E)�t0�%��o��k5�8��y|(�{�<��I@�w
�-X�wun�������X�c3�e�[�~��蚮��� �u�����`�ξI�d6�?)楝����@kp�Rz��Z9��a���p�n=���u�m�I�<��|J�<�fėg_��{��F���&h�=�hp�L�.�6i1�d�%$�X��_8���k^,��ټ��4wp��#�D�R�~#ZkK_Sӯ�T�!jx�@��x���N�n�j���7���OF%Y��ɛ}�����n��Y�I�z��/;tm~����ͳ��̻��:=�҅�j�oI�� J�L;$7Bc�$�"9� ����ePF���������/�i/K��x��}��ॷ��yn�,t�H�BEb��%^d�m+Ux�6�$��>Il�>㳑�`d�ʁ���Ep˩���v������`Lm�Mf�P��p�|_�/ ���\ܓ��a��jcjƼ�!tK:�,vh^Ŷ�f��E��렬-<�yp⣐m��˙�C�3ߟ��yK��лe��������c��릿Y�=@)�;����E��N��'��^��h�)�g�~#�Ʉ�yG����u�0�^i�؃���ޟ��y�zA�YS�����S!�ao�M��"g�`���P��= ��2?��o�f�f'[�m_!/a�T!>�@�Ύ�y���d�O!���yq��Tw;�W�Z�my���������%�E�ƍ��;V���^�I[^_�{��7�"�4?��K���͇5��W1.]�[�x����0�##F� <{������i[>�v2��G�8�jp%����+��L����?� ��\�>���W%owT�j���/���[x@��h��(�X��J���|^�_�P��%g���(���3��?����"��`^��~��:�� x��ڌ�}�}��ʁ�+x���A����ὭÈD��b�4�[�<��e_l��ح��^u�oc�a,�3�u�N����	�$~�XO����!/ю!��
��x_,P��.����Vrb]+&u��)�Iv�/�\���E����rd�A�L����ѕo�w}�3=Q�44���dU��F�
�8/b-��$�<��p��[�����d�=������9��^�� �n�)�R��(�Aޤ)A.o�8`v��|q�fq��{[�D���$F������Xc��O���e��߁�F-(�G}-(��	�-���hM�{]�����Q���F��4@G)�2��*?�(,��ur��Ҁq��h^�&����+~wk48uރB��{�|x5
�0�6D�݀<�Z���){�oY��DW4����6p�{z�^�y"������*EVkw��/Qhƥ9\H���xx5ۅz�.���3L��r�ǝ���1
��n	����:�n�Z])��������<��X��Xq���!͉I/����R]�mGA۠�1�j�^�	#=e��Ս���>�I��8e鰵�b����L�2���<����R��dHJ�.�^�Kʐ�/D�e��8V��x�8�j<��{q�����<�/�E��T��I}�A?���YE}���G&�ߴ".�DW1��4+�dm�>��+��ÚJ�}csm�ሂ2�� ����r���$�"�� (�
���Ƞ�AeN2�`��9B�H		����>�{�}�{�����^��?ػ���Uk�֯*U��!�K�|�>���u�O|����^������Z��OE�8&-q�g����`�$/��UJj�L��I��X���/r��
�3�Cف�[ �6�m�F�.J�(P*�;�Y��h�R5�W�\">p"���-�0MEɜ"������K��݊����R�1����&��S[s�#w�GB��w�z��p�߶�ZYZ(y��q�q�8�eu��9Y`1�w����p2Q��`C#""���1����o�#>ǳ�D��Rֳ�9l���r;�*P9� q:4�i˥L������5%��@![�}9�&����Xÿ���}Lx����<Hv�)_N���6N�7�(��^ڑM�.ܵ��뉫dĤ��ޏ���q�<9���=��)��Q��&��K*�|#�i�S�c����%����_�R��9�k��M���Y���礪�+L�� D��7��+ֱx�s���%�������	�m	7Ʈ�~@^����D�$!����0��7%�3*"܌�����Y� .�a����~E�M��`^L�G7�� ���)ϛ&(��t��|{�1�#[�,�6��4e�����z*���lI�����V֚�=��V��
�Z���K@E�u	X@�oR�&[Q7�(�V���+u�P�5�<]�����J��=�Z}턆5d������9r6����b{t�AM_;�߿��i��V�Ujxyɸ�S������ֻ������w����>�I�AG�����;l���$��`�)0b�ʘ��ϗ�T�M��2T���@��W�p���D�]T'�'�T�}����M]V�|�*L�^oj��$�Q��=��7�U�1�r�=���!�����ʈ�2��[����I�'Na���-��Ũ���٤xg�z�����g��U�7o>��Rf��j�Eǃֶ�k�y�'E���`���/_'R$��f�A8(XhX�L��Vg[� ]��%/�Lꥬ̮�T��7x禍�i�/��b��~U}���0p�&'~����q�Ĥ$�TI����@�c �c���P�_*��3���B��*vtx��X�WK����b��a�j]z�������vk�u�2��yy�k�I[ 9ΧW0�`1G{=巽�o�K�.��Z-j��U��`*�`�*ʠ�ƛ�yܰ:i %����L���]:�%�ɐ��J?
S�E	��f����,�l��M�'��7e�Ol���>m���)l������N�eׯ�N��W�Lкk�ޜ�?}�����4��Ջ����tf��!5~Csssg�����2����@p��7o�H�D*�n����B����|�1��=�o5�I�M����%���QdT�ߺ�`$��볘��$)�> �׺�q�+K֋�L���*L�ș�Q���,�[a�p?zt�Mxa�J_���6�`��m:�P���"�A���Q���{�/��L�J~�?pa��5�s?�A-���G�'MB�`��(�r���`=�C�%�I��~�q}���I��58�����In���
��I�=��c�2�;66V;C:�箏~�FV	��E��*/\�/�h�(!����	��N���( ��R�^h8m�V�Zu5ֻ���?����=Xuwa��z}o���q����ʻ3�X	�FN6�N�q�n��(����3��*��'G))'??M��7ٞ�:b�J��������\�n�u��Q�Ԕ$K����+�-/�RR����sM�� t)m�`շ�r��įC;�S����K�%�g�'=�OYs*P�U�o�Ye�n�cw��s*	@kq������G
��V�I�A�k�wDM��%��0�B�ׄu۶��:���!�#:��J�_���>Nqʦ�I\�'>H^���#�7&���t{�>����c,���MMMSA����=����f��x�Q�%����P�Z��2B%��e����6#�l�hnz�p]:p�����s�-^'�%�g̸|e�v�R&�`�t����z�� 6 �o>�Z�����ܻ _I]�5�z~q	>�C"߮l(}F��v��{%�M>Y���= �W^�t~r )^%7�֑/	�}����m��b08{�=��>������Ѫ)�:8���*�D��Dݵ:	��'���_�I�|q�̊i��q�1��$Z���� %�D���5���lRMpP�	Z�_�	
{�}gǴD4�l1�=�3�(U`��OB����S�,e�4�T��	�jev�y�����O~|���(��c�5��.�S���#p2<�s1�[�!ǎ���D�� ��~�[�!sC?K���Џ1��Y����2�E1�PU�����`" -#�]?���a��G�ېW�� E���7�_����L�� )FE�m���V�޸�)��X�:EC,�߃-���ץA'���8�4F2*Q(˴|�?��#�M4�x��|Q&zௌ�P�N�Q��~����ba--n�ys'��*}	�|��ězg����vY	�(�@'�1���eC�����8/�j .�q9�������ݤ�AIh�(��(WG0杳�Z�A�g/����.�d	�$��1�.��ԡz��@�s2�`ʳ/*�5���V;fQ~�:Z�"��{����kP�� V�ea��a�ꞿ�̿����~����Q#ӡ��򺓐b)p`�`�P�fЂl8�ֱCPV9G(���hM�eX�[@T�G8ȫB/�A�Yd���}������o4fL���4&Y�f47x�ɑb���H��A|��(˳�f���{����luEb��(�b��*�ΏP��
��=CN,����+���b��RF�+ �d�I�i�r��q1�x�4gQog���{��S�l�'�;��8<,&.}��4P&�S�.w������I�X'��ʼt�-?
Y�ܯa�?���^.b�F`b�;qaf �o=
)�x�a	j�`��� ���5�����_�	�3���u�2��SR���L������/KY�����ԪP�\�P\D[�@�{���;?�׈l��������W �zc� �جm��2�kGA�g�wy~tkG�ڭ�G�[�Y���.q�r��zv�a�:��-�:J^����On��{��n��8u�Q�a�����L�����%��V5��ѡ��/v�Y^��"hSa�Y�#�x�e�g��D.K��/�����	��Ē(Ŭ��&�Θp�s�/JpM���Ж�^�ho���R�sGǑ'�!�A�����#�=J�����c�OR}e����+��ݹ��F#Z��%g�����wkoƄ7ekdtU��q�2�*����9qC���N�M��@0u����ʯs����JY���=�B}[w���??w$ԧ?�S�iA���y;�0�����bL}�>��+K�>󄹹��%��O��<0�Z��)��~�#���dۚ��V`��R{�����jT�za>��n���l�n�-��Ź��=t��[ny���|j!�?\g�v9u���ߤ�z��V�\h��%�ۻ�љ����i_)n���^��]˧��۝���l7 ��}"_��t��7�]����mK�8P��60'S �eೲ<و�#��(!��3��u]�Yn�l�v;��U�S�"q�N�[���NKd�(P:ҥ�����n�{�\���>B�����۟5�Bޤ�+��E!������'[����y�e�O͕�,M�;Yj�GFa�vlp�U\t�(S_0�r�.r�b/\_�\i5�ф�§ϫ�''a�~x�;�E�͠���龧gTc��t����с�n��B��2���oܫy&m���#���4����z�y�W�����s�����x�@���<x��R��y��CJ�	��s^�h,��P�%���sQ[���&��G�ܡL�*tV��ǫ���ݚ�:d`�~���ߒ��d�6l�Y��L%<��������v>^��������|�~�ͱ	xw_�����D�IYz0����X�=ٷgg+)�{M�P�)�qL��A{���Dn�*���=/�caFH��J��~Xٴ�����ħ#�"~ﮪƾ�%%j��[�@'`�^����D2^��d[c��@Ѽf�e��SS�������`�n)�:&�[͹������XI��҃���vS�^�g�� BH�����j]�Ε�N�N�c~t��^E�R(O]�^�΋��G���,7@�t7��1�"��}Q�j��z����5�Qx��$��Tp�K^ań��J0��_�'ʑ~�A�j�8N�F�z�d��e�G�y�ȧ����HǌS*OZ�;�W\������"�vnTۥ�f1������=�� ܋��c�V��S�(-�2Y1�%a�/Mt���jl�JĘ?�|���J
S�e\3y�Q�,�TQ��K���@jq�=�����]��&v䒾����鞯�������8v}��P�[U�ߣ(�=">k��f�߂Ѫ2�͝����N������ݮrB`�/1Һϝ`��w���	�(K��5���h!����β�X�D�5φ#�푫�r�3Γ����>S��"
�P����`�n�[XJ�d�ݍ�Q�+�	>�8NF9�|��H�qMۅBX�:?�D����%U�V����V�Ǖ��T���Ow.��x�\�����-o"��ӎ��Np�"��h�/�mz�a�+��Ƙy�f9	��o0WR����c0�	BwV�$�]���V�*��m�=��~���|s�j�/aV���+�h�͂�R�w���w"���,�|�Z*�c������\K����Fy��yZ@1����]6GU)ڨ�!-�#�Մ/"��������?�����ZU�ܞk�P�?�hmח%�TN���7��1J��/,,��'⸾�KK{�!�/�vZb�����5s�@�W� �������C������g��w}�ϝ?O���IY��J�����/�,?wH�ym����{B��#�[δ�d��kM3�gΕ+W��xw}~��d�G())��\5��֋pL���p*;��9��Ɯ�,�7�Y���&C�lt��p���s]�X/��H�rS.�a����%���$	���@uD��T|5����gn��OC�׎U�jp�Oݭ�΂;D"����%zy��6���z}'���"l0�n�^���|L��	��o���R�܉΂�߱E�-�}�l��3G$�;�w{�݀��c[��K��b���ӥr���p��Oa%u����'{RRR�	�$��mwf�B��<�P���Ca�����au
���Ȑ�A�ڋ�i|f�P�ѵ�Ę����|����H��T@��E�{��jk;̽��E�D/R��H�b�xOk�w�|81ϋZD�Aj�� ѣ=7\_O�L�=�'�)l<?�wTC\N�:r�1��7�`{��ɓ'�[�����E���f��3�-[���bC�k�����	&�(�|ľ�3��O�$IzQZJ�@�-��Oii���!D$��W�G�����a��偺:RC����OpZ	 7�ؠ��H�Ș�؊O�=�~���	��(���"�j
�=m��|���+�
�϶�M"��	߁�d��$	)f��������S�q���i\�~��-�`�r��y��ڍ����].L���r�(k{{�&X;�#��`��-u�0r�X0(�N��������e�P�(����lœuTu��oAh�R�����f]z�L���$� ZG���U#�kݽ��=>=�l�5�L���f��/���D566�h��ބ�g"Q���=����ݣ��ޚ�����EN���jp�77���J���`�+a�@�m�3�������G���Eq���d5k��UH�<H��s�v6��|�S�-s�w�ퟥ:Gͮq�дLX+ru<^�#m|��s�	��75&*��;��[�=�o�kD�����ve�$�]ײ f���9�6)�U�^��e��U����Il�>������t$]ۣ3�bb%�Z"k&�?�2�����g��X*A7�	'D9��

bY_���)Y���%�� Yx_A|!��;�� !GwSJ����������D�Ae�e��@
�:9C?�)�ޖ��������.]�e�p�,,,h���َ�@��Q�h[*p>7����-�b{�g���Ucŉ�/kdtv��1���a(*��PfFZu�R}���A�d闓����U���!�=ؙ��E���v��3��a��q�0#�Y����?�$	v���g7h�ٓ�D�5|>_` ��d1&'��}m����H$R���Ç �|��
''';�-�7��F�^��K�Iutuu�2��L]`l�O����eH���G���ˋVy�zb����W���k
��O���Tuh�k��i����]y1r��g�s�E�JIH���)��?�jS5�Z%��M�g�52$��;�o�E*4�����Rw�rLLL� 4Wfz;::bhA�,�1Mob^��[����?�ژ�pSo	*zC(�Z�kq����@=Ka�ь4=�2�R�ޗۊ�o��	
rd��ױx
�z�9⼟*R+�Zx)q���o���}���I���PK   �sX�X�޿� X /   images/97f4dc10-5048-4749-8251-75563a783bed.png��XSi�?��NpG���У8#2*   �A�� V�"EB=2�D���4g��� ���(���PT-�HH��9)8��������{�^��y�]~�~���	�$�Ӳe˄��5�X�l��e�~�Z������[A��o��Ǽ�-�6���|u��]˖�_��`�!���S�����~�?����������*��,)y8|��������*�ݜ3�~�$��-Ş���Z�1��������ǟ�?�۷^|���?k:zy������p߯5�!OSqa��}7~���g���ԧFA��Fr�$������J�`��Ê�(1������5��}���6��5��.�I��޽�{���I�-c=�+���eBJ����UY�E�`Z4/8�Y�Ú�2di{ ��E8L^�:M��c�a�w����5���6��娿�;k��4x�챲i��L��I����d???��W�yU�5��4���#��P������-G��>��iZ��)��fbL����������*�����xB�;":���ס�ޖ����ђ�>(�upۡ��y�z�$���'�L_F]Q�a�B+�Ɵ⿩����h=�
�*@�Te���Bb-J����9�K(��X���7.�n7|�~%�C�q"�(';��i����D�D��M�;|y�e�e�ź����Y#^^^aC��>�.&T��7����/<j��z��n�,"�JA�n�"���\�QỊ=�W�$/��!���F�o(�(⍗	���R����	�7��zܹ�����(��΀�*(��(�j[n�<��:n�-�&�m�����k#q�أq޽~�:�����s��`!R�����1�伛�|vU��2�mre����������֢����7eoL)�(����2P����"������J��� p8z<$|>����ў�	�~�g"�#��E�~����u������PhC����C~8�\�|ty/T�g��Z)�w��2�R�>z]v�|j��@4�=��s��y�>>���xNCJW
�7�Z(y���j���]�[2$�F���v���9�CVVYv$vq��?X��E�DQv��<��"g�X��
��]syvM]3N<����J��8�h�u���u�/�<[z�N��.4�����?)IHJ
��֤

�{���6צ���e�۽_�Щ8T6X����W���D�����/���C��e�@*pj�V��p�
n�A�|���b�R��|o�>���SF��(�$H0f�Q�O�~�UӔVE��\To��ۺ�?e���o[a����N3Io��=�����֠��Z�~qX��333ML�R}��p��b[�:�Z����uSeU�.��E+�2,�-��y��,U�VVw��EI_<���(��v\Iߓ�2t�?��p����VV�5�@�쪶e�P� ����%�,J��Tp������/����:#��{jb���ie�����븥�&~�S�u�$&�2JR]�����e�;d����� ��D�j�˲2�8`�u��x��w��/=��}�����yp\]S}�R5�"vΘ�����]�����W�C{n�����U��0�n_�v~U��9;UŶ������Bfq�6������,,��f-�Y�����)1�ƔN��kp��QX(�:��VM���/-e�S��<�+�z�e�m�X��)7�sq��p�����2�Gv�ǜ���kpJgLHJJ*6�{H`Lr	�I��5�@ߗH�b1f�":՗8	e��7z/�A&+B�r��?�	�]��V]]�Tߡ�3O%�[���H.�K�ђ�8O��kmmm����7��,�z��_��L6�̵��$O�:�Y1˺�g��Ɓm�e��7�G��WyU�vO� �V���b�PVA�5���������Pc���݌�`ۆ<���wK�9�x�H���1��A�O�F�'Ux,I�X���S������^31)*���b���Lў
��A�] H"� K���ݜ��_�"���T45��
n6�yX>l�m��c��gف_eC����?���ߧ�˦�4�\䣋φ�F'�aM"a�9H�p�0%��cM�!���d>���"���@`�?�������;�O.,��^S��h�X�u��M��L�g"gvbKe��B��VVv1<��;-ν]��[�E�u��$P��N����Ҿ�	���|`�:�,Vx΅ʼcϢ#����ۯ��̵��ǉ���'����NLw���'�kʆ�����T}��ֵ���vivj|@/;�>�ni���^��R;�;�����"��=H-6տQY*�C~~~2&�!� ����A�I�H�<����$o��*��n��ί/!������qS�wvհ6��YS=C�wSW=���3����ح��9t���ŶX�iY ���{	�4��.|��K_-�a���i	

:W&�$3���5l'�*�q@�ط8�U�}֔$��[=�wM��0�Mڳd��+�:����,u+�����W��������j]�N��i��iΓ��Ա���
�R�3�P�m����'و��	��1��Xn+y��@:�H�*ٶ����E�h,��w����-���?LzK�#����r�\l}s|=�˻�>je5�r����^799�2N�e��?�̰�+���i�*V�Cq��o^_}u7&d�ޚ���d��WK3�������׻�̫�"xKSv@�<���k����e���&_�ׅ���j\
7Չy�@-G{���N��-)on�kh����渿 ���W�S���/�{�M�EO�z��ژ��ka6�ӈDF�1E�R�;�v�u#�e^��Ǜ�z�i��-� ���Jb�)))MF/���,jaH�������7�m�m���sj�!�F*�D)�$�0��+�*��C��w��x�]顱5���X����.r%_2���	d���]<O���[��tp���k��	����97~t�����r}ٮ�I��L$��{@B�!+�OS���&>���sj�=��j��@'<0��]>��oHg�x]�`�����A��8��>�:�sj+��*T痞����y�pu���/��#l,�A�s����O���Jkc��ۛH�eّ܅zł�-5��r�(C��i�w�9$����]��ɑ˗B�I$�2����Ⴜ�6���?}�>5fԴ���L'�T�=o�T�lllL�g�"��Y�-ލ��1�9�Tk޶�W	�@y�^is}}}]_TU��$_75�A����_��!���r͈=5ک�ɠ���/"*�~�h�=5��*C�pm���L$!(��h>��Zp��"r�pM��^(����C��-m�J<�=S�9��@�M ��9S�����~�ja�����Љt���Y4K `�=���0?Ч����{��t�/��ч�\�ӊ!<��:���������ArhE��]�`�� ʈ�����2�\���9BA+8��Г�o��h��o���t�v�k	�C�z�nGu
��MM���гyKV�gV���ޟ�/���;����gds.	7�N��;��'G���l��8E�����k�WI���|�,ݹ�}bLs�m[,"8_ XIIa0�ȋOq^���⧵��D�b+�G�����D���9�;��_�*�L^_^axJ�NyA��͆5@{_U�V�7��dl�=�]e?�(n��>��TLC��[y7��Ӈ�F@^��(���'����u	����� n��}/vJ�V���x��ěr�ƶܔO�t3#�Z���0����H�P���I[��#)�BR.�y:;�<(��qJ{|�����\��Z[{�9�}0v���p��]ޖц^���eaf��� �=A��������ǿ��+�-�u�V�~eԞ����4�p+�F����С�i��čC2�!�Bܧ��9��A�~x��7��+V��F5r�m�0m�P{�$$%�᪯��(:۸]e�N�D��2*���q���:Wc>�uW���E�ОP;�b�Y��I�j�z��/���{���K"�6hZa.I���5^A�����*0�z��_s$+��3�g�l,����5�s���4p�g�k�t;������sq���a��=�7�U��/w�����ޥqLL���vYv�@Y����c�����C����͚L0�fh��\�G���F���Vt�it5W��Z`�N����F��4����_	�&�Ї��`����ǌϠ��tP�>du+�5c��Ä�+�C�7
j	'�����$�}�t`y���W9i��"�&hZ!��4��4uw7���P�Y�K��#������;`<�檗�PB$�C�)�ڕL@6��$����VW)�L%GgA���D9IX��`D�c ����M{�Z�����ٹ�r��<s��@��. ��q'����z|�v�p��ͽy��s056	� � �6yZ�S�����
��}p��7�ڡ�e{�ɳz�]�ا�^g8E�J�#|b�ik�V�4Yd���q�^�h�?����R�=�$�����3����j�+�#�f���94��{��w�f�s�-dv)��G���sv@a���#��,'�C���W����4��X|()�H�-N�%S��ء��L4�h��qy*���r_e}���z	U�X�\M�ZA5�eJ��ۤ�v�>�ۥK/�-��>�eW�SR�u9r���R�پ��C�#(�[Y�3�Wm�:�>���נ�.�@���
�}|��(GWY�w/�v�75�:Ϙ�AГ7ݼ���aTȕJ�~�t"p�kD��̓��e{�	���N�F�K{Y���D���X���X����-��8��QDEIJd�)o{�۵İ1Vyx�v?5�k �֢�e@kx�������a�y��C��PF��h�����yP�}A���囸�����1i�D�C��0����h-{�s<v�g����LH�/=��q�ww�u�w$q�^Ԅ+kl�[���v��Q��0~��N�Qǅ���pD���-6�V�T9[F�����Rm�=A��^��a.h��{�Q�7�m?W/�������G��u�����tp��SI�F^�-�ۙ^e���	���<�|&矹��!֐���A������H�[�C��"o�k�EVw���<9���������w�����|rL�k$N�i��NK��%YS�j[t�	���Y�ų�>�"����*%��NW��k	�>��*(L��pǣ�����ڽ��i��������-T���*�q�U��T�DeB_�yKn�Ӌ��T$Z0��{�?�aR�G�K�iմ���ɒ0�/(�������{j�9?z�H^Pn+)������嬬vD�� =+d=�������pw��ҵ�ť�Mi� �A>�q hH��̶�bE�=Pb��K��æ=���e�Gӝ܇'��.��}���*�$�������%�S��o�J�rv諫�_���[��󾚉ԴX��k�WCVVj�r_��5�ni�#��0glP6��^S�Sg�Q�B��u�#J�j���B7�{!�b?��j��k�n���	���M�3 z'�jj�um]eT�J���4���x$��@�6��Q�=`��)��|�q�˄�U21D�M�?�o��mE���B��2[�2L��|X0q)�Rc�����9q�<yr)��h��A�/h��!1*��]��k�F|4���Y5��!Q���/<ZJ�����i��u� �s�r�c0x�о� �07U��7����N�I� G^��r���L����txXnk��0�B{�
Oh�G�ʘ��.�P����T��N����I��B��v[�r�z?��S��Έ�\�v�L����T�1%��D�r�zi�h~��#3����Ez����#/+Wr�d�5��7�9��AlJ/�?�=�����x���l:��[�(��e���&��@����\��bS�3��+������Q�uh��KG������۝:Po��������ӣ�;��򚩦�?�7q/�}is���� ��ݣ�YbAx{;N)�q�]Y��5&.��ӿ��W}��%��U��(�Wt^���|��U�A:s%l.�#�5!�ۨ�!��}�`V�x6|��J�5��H���-O`���9?� ͈	M��qiJQ�հ'��mܯr֤�d���U�#tK��HWY�^�>ຢKLS@�5�(��ɛ^��ټ��DO �rז!%X��&݉a�8;1��{%����!�L�ꄫ��b7<l���A_�Zo(�D��r�*B�vn��p�-��˺�/{ƣ鼑�Ɣ�ȇ- ҙ{eG�
qD�G�#�Tzr�#���V��I;���#]�`}O>��I�"��:�q�j���N��z�S�j*ԋV~]�&eXZ����^XL:�߃�4r.JbVe@��n9Z9�6�;�}�D�jcϢ4�͎�"?UTT���8}������u��J��������n��XhƛzOA E;�©Yn;�=u�7J9H#?mf��s��8���r��6h+;`��	�	I�V��Q�!ԭŷꎌ�'.r�M ��'a Â\�r�~��+�<k�����.W�ųs��6�����egMWG� )צ6���{�PO�~WA��TR+�,�X6�lc5��liL�L�nhՌ�#��R�ݟw����c]�W���9���Cz�!�:a\�H�t�lRox�,�TJB"�(�5���6�QyW��he�f�Fk"x5��D<ܒ�(>7-/t�+=��(���c�����O�f����Hg�b[���B��q����5Tc�n�q)�M��]�W�v�����kx���i�S�:s��*���STR�2���[���_5����Ҫ��Z�e��p�p��q$a��tJ�Vz�_���9ʸ�~H��ΥkT�{Щ�G"9��T��M���{p���pPfhʺݗF�ר¼�c��[L��f�3��;|5O��k�Q�����Z})G{�V.SG��VN�ǝn�>p����׸�
,��"0��[Z�o�+ߠ��Y��9��>��j�T�2W�><f��:]�"
*2E�8 ���T@�H	t� ��K�����\oK�Z�6�0&Ƀ��~I�zQh����!L�P�Pf�mS�#�5Q���E�j�A3�
��Q� ƾD�#)����Z >R�p5�缌��%�儹=AIPĐ¹����&k�v�a�1^,�����/�.��*�e��L��Uʘ"�*V�~�2�6iN�f����9�BF����B��^'Qn�a:5��_��X�_ᗢ�㑾����1&�l��_^�ΥcS�}�s��>	4k�h� ����L�D$*z>9*ſHl�3��^�5���謬�I��N�6q!Ժ�����*��٘����n�怢Ν����[r�"}���F�q��6�=�}��ǛQɘz����(Bz*�TP��{�\a��moz��'�o�'W��<�2Gm��3`�ep�`o`����5��#�W� %�ՋnP!�{�ө;o��ΚKY���6;r)�%�}B<R/�H�"u��E�yF�#rj,��t80��V��jI��v$�l�9������L��ܴ��v�U��P�|�]���RkvR�6�ر'>�8��Ɠo	�B�UB�_��ƅ>u�b�a���s\	�+����4��x���M6�ɡ�O�������n�Q�����-oXӅ������q������m��{˧���^�	Л�GR�ogo�e���K�:QfX�ǜ�`�9�(y�ѩ�H �y~�@�\��L�o2�?��U�d�c��h��@/�!���[��m�Uƿ��^�V��vo ��K��VH��GO�@,�������"m��eq�=pd�T�kr�7��%cy����c ��|'�^toP�a�f�P'I�K+�,TI油�ޠ�6H��Q���b�a�w�>��Cff&�t�#G���Zpg�ȷ�q+%X.u�fK�p�*���B���P
�/�՞��&���̀پu�~�{�[��)��9�M^�5��hJ��e��������2��0H�ݎ��������O�Á���e�7Y� e1�+�6�CWAa�g��-���@5�{Ιs��#E%�:����}s���@���_X
�L`��QM��yj	��*f�H��������3��B��j��\{�����c�-�����%�ﮂZ�(�Ŏf����ݴj�E"����H~|F�3 ���;b�N=٬{zz�B}e�n��ͺ��Y(��y�hLU.+\Y�&�ȳr��j-�����H;��ņBg�_�̹�&�&(6 [���m��q�/oY�V<�Й)��|�-9$4�Yg��0^L��061�7��y <%%P��|�ʊF.�\��?@x���@�Y����R1��y���V����u�S.�P_xhle3���R�S����MɜqJ�����S� �(DY3�em��=�e�/r�"q v]� ��!�YY-nH�lJX.�?[?DBF�I�
�($��FЋu�yi�U�텐y?HdV5�	K��S�R�7�()�t%��e�R}�x!
�ųfHf�!$���-�d�k{0�YL�o�����x�k��4��0�eOɠI��Di�$��Z��0D�J��0�~|J{J=�+�#�F��y�ߋ?�BI��#��]KY�B���f�YYY�H֘Wcx��m���1���X��b>/��������OJ�j�RWN�:���Ӽs�\�<����)F�B֫�DK���?�>x�gϓі'{�]x�Z��p�jf�4��F��u��y�Se*p3&'�vJތ���m!�~�o���q�5-�з�Z|�j㞲��C��%��.ő�Dbo!�	�h��{m$^�G��E�r��6�@i�&:̨�a���������<���ʻ�6omeEJf�U����M�[�4�ZDWq�3Jg*��(~�r�RI�w���G�p��"�?*��L/3����O������#��B���j�ƞ���N�Q��j?��M�WXG�CP��/c��hL�pϒ�9z��y�{\E�Àt[n�C��v�FH8�qu!;r�nm����+�#��(� �[�HW�[|E��$�(j���hB����<��b`8�sJX��т.7�_'9%�v�j��?��i�;�X�<�R�[4%����u1h|,�
��2�#�7������V��i%��)�������fke��wD���F|�� ����T}�!��rl�Z
S�������ˆ�Ȳ������&/� �mu���r���~�v
�[�}��)oy�v1��]VV�Y�a��6�y���(��D"v��h�\��$�^�N���>U{jHPA�vb�^C��o����5�ƺ�����,V��
�ӓ�s��F�b~��.�@�s�u\5�rR������:�9�[�.�j%����Vh�'�7;���uE�J�rF�O˭�ڎl�"�VU�r�t�*5?�x�kH�8*�}@�L�SZZZ�dM��b�-q�[d��@�u�kOv�i(F.�y����ˣ��� ��A�E��������\�p�X��0Ҟ���1zRh���z�M��/8}��=�E�d�a�UְF�48�2B�˯t:���]L��"t�l{+���$�7b깂/�{l��ƪm�{��(�p?�i�xw�b���'��Url����B-f��5�{�q=��<Cg�p�@r7����&��1��K����F'��e���x�[�3�s�D";(J'�5�{��[�A���0Q���Ҵ\�n3�3�B�W8rF���4w���̍QO��]	�{i�gNWW�!��.���=e7Gf4C��4s�S��
�J�$2�;1g@�O���d�6s Z���Q31���h��&������� � x�7��(�֕qoҕq�pj�{���	~�l{d�,]�.�������|0�� ��H�;� ��S�<�[~7/az���Y-��3�� �3b[��K�ӓW�5� t���Z���ꀸ2α�C#b�i�U��,&�&�6�ϓ{�@���8.�-�@:��DR�Z�JԪݺv���g�(�Hg�l�Vm�\���t�wqY#���ݗe��W?�G�j-�=ۨ��|V�Q���
���Ӹ��l�,\��X�v�n�ch��5Kg{ֽ�FV����7z�]�`�e"��� ���4��~���,��[:��ˮ�N:�s����t4�|TT�QU�o,�XJ���l <|Ժ�z����N�B
S���?�G #^u�UM���q��a7%;�tGm�t�w���0ƹ�>y/��EΔ�d��T1��� �!���R"��N� Ot��&�����δb�6�*J�8��be�2ȱ:^�y���	�
��ĭ�!�Wp v��ƈ���t�E����N�8V��V�Y�~6�j��8�r�I���S%ճn]iԷRҜ=)ő�]���B��ֵ"BZ���	8o�9��r�TH����k��2�Vd>v隭ڣ��B�;X�%[���N5Ơ��d�)����ؓq��b�W������vsOcc��Ɓ��M�a�?�~2ⶸ}�[T	^����(b��Ʋ[��CH�yH@��/k�T+��2���8�k��,�o�C��e���
sZ\e������]�Ya �1�n撩��~.w����aާ�n�:��^�="Rܚ����[��� �����G�9��fW�§�\��ZR=@��QowN��A��6iQ�ˈD�<q �1���]�I#���BE�q��<�߹s6p�T��m����fҁb��ڈȇ4�#�`�>B�E"v3�i/���U����
�;G���ުRYy��+�	��K,_yOk�'� ;��g-q�'д��P��o|<K�J|�NE�?9�gJқ8C���O�-Ҽ�C���Y?HH�9��Tm�?�g�i)�>WJ��%)�4X��jM�-����A~D��X��kU�i�`��U`\�Yd�"e�1�)Q5��~�8��{ʐ{��~}\�^������ʊ���9~�����[QNy�`]+e��[Á�s����Db��l�m��-Q��'���Ra�N�J'�6��dg�z�32�SC5��8��9�V�S)����RN��[(_:�%���P[�����d.�O�"` �t�@}�'�K�� ��"�V�C�%��4a?�ݲT�%��b� =W�	��8m1�aT��$�7�?��F���<����
��?�366VD$�L��ۗ?zQ*�4���x��[���/B�I�/@�������Z�S��X�d�4�.�8�(����^ڣ�z�+���~�ͭU�6�D�ş��cu� x�,�W�����܊��p/tT{@�M�S{��|ZK�[�YYE���'hZ��'"�Z'��!�O&�����.��ar�4���my�L'$�n�;��pwOϭ��>��ꅔ<�"C���#eq���*c���R�=B�k H���εV�����MN�y��U��ؽ����z��pf�Ν�M��͓k�@������a��+������}Vݟ�Zx���tk�Cg"deq�@Hw?@-�V����_�(B��3#~�I�!}j*y߼�{�60͒�M�  v"*�5�6?���,�,��W�͟<A;!�q�1�BZ��uh�5�E�Yo��ʭK9��F5ak����Z�Tgr��������lp��^�<��̳���%�6~�O��f�{N2�+u{�1�Wp#��:�<� x�F¿~�D�r-����ʳ��C�tR{,ә�%��k�����0n���EWË�� �����9q\�=HC�Z���.�����OS�]hZ>a. �iT��D�J}���sR��N�{w��K����Nzz6��g�����f�H#�)��z:DDI:�=Bδ��dA�9��N��ۗ�~��	������fk�2H�UM�e�GKj��s$)�E��l��L6A��,�+���SI$�ӧO*���Y��|"�5
aՆ
��Bv1z�cI��x��<��I\&�����Y����u"�������s6�Ŵ���x*}�n�􄧌sq�C�P|6��>�G�9ۗy{��cǉ����{j��&7�E��%�[A��l�c�Q���t��!�j8H�Z4���QH$2�,�
�@���U�Eܓ��
%B��7�e\���ZKMծ�G�p��kT���{�i���`]�$"&9�{��R�W>��"���3��Δ���C ;oBZͯ����z�qNSu�y���쐈�G�_�췺A��1?nmi����b�{MH�n��H�ͷ��kT� �^7YO�__;�c\��;6�F!wl�q�y�i��"N�s#>���T*$��9��?~+�LT�ftu�JH�8L�ҥsM�B�":1N��H�n`�<��c;|կ�
w��C�7���]������ ����;���(A���ҽpKu��Q��'b�T���_=Z�[�n����k:^�׊�A��B�$J]��9x	s
q���G�C$�4�k�Y�Xl��K	(8F�(�5�<|��",�A��)���˗
���Aj$���7�˪G�f"���=r�Z����ٗ�܆���Sk#/����`r�g'��e+V��7X�.�EI��;z7,O�B\j�ȴ:5�U:�D"��i��!H-Erj�m�g-l���G���#I�n_ �ۧ�h0���zQ>F���eI�(D�_�L���v������=�<iS��	��rf��S�5V��|5y�
��`�q���=О_]��w �I�9%ȟȐFq����'�?	4��Y$���`�e�������D"�e(	w���I�S2���c�i&ޮ��ST�d�2�).�«�V���qWF�qxXZ6hÅ'��ض��*���Fy�3�����8qQz-�'%>�)5�j�a|�����"����y^�q ^� ̅��(�SH����rщD�{�ⳝ���J�����m�c6�v�al��Kp�-���xu���C�pG��θ	���[��D*�>�9�{�P"�P"�7�\�
^9�A��ZE"�,^�2vg� n�;{[T������ؓ��D�T��n�����Rx�?�;�;g�IHv������4��{�v�
��t��p����zM���{j�n �v�,���n�yc�B����2�W�l���a??uc�-���J]v��0��8�Gm��f��6I��v®�]�er��SO&bTm��{��5�����Fg�R��
��oq>��jGp�4��1n�z2�� ��2��k�=nQXX��P��}�{�^�Su�Ĝ�f$u==68)���˸dB�)h(�kk�ed߹�kH��y���LH��O �1Y�fX����ӽڰN�`�
�y��<�]qԪ-�\�qV\G�Z#����N�Y\5�0��NF`���@�`o�u����R�E�pa)�dPB��h~֥a�R��Ȗ[S����a�d�{�p��ަz��������j/��?ɘ�X��k��[gk�A�YL�6�ԉd���	�⮈�D8v�R�vT�~�iʒ׆)o�6�wbN���{;��ԛ~¨�������Si���0�h"�~|�ڴ�"����L�F�aЎ�k7x�F%r��ƙѾ�?p���ØL�0�0w��Vz�b�0��r`����nt����;�9�Ĩ�����1RA�� ����)%B1r�w�Q]c�f 7��U��*��T�E*������l5d���0��|"iT	=-k$�_K=ޔ�%-�˅��=5���u�_�7_<�3��	�S,��u��К�vg�{���BV�!Z$C�v��$[��76v��k�JE>ڠ�m<�������4���o6�����`$���G4Yc�-N��l'S��c����5h;a�:�0A�z|�9�ɣ<p � �����)��e��:Fx}�#/�I�8��$b�n�����$o���}�c
q8Be�y'R,;�mR@$R�� ���� �_��[�B�&��u�����@E���ŗ��(5\���Q���$糪���rpʺ8�mܭ[��pN�$I#��z�CS�5�0�z���I��v�?����ɾkX�w��g�� �ʦ�$�&7��kx�k.������5�;�dy(J�`�x��k��T1��3~���0�ږ�
ؖh����z�3wA�܏�b�l���7[/�Ct]�Ꮢ��y�>Ңj�袿�)A67%��P��0XH���3�\YY�%��]GU���"���Nٹ��F�����Ձ�G4�����^�F��A�]�)!�CM��^�@ʼ5�m��8 ��E3bG����2�>��2f���t0���ΡiS����Z|hG����M�Y+��; Ѕ]dVoR�c�����M����q%o���̇�LV�X�A����2�_mB'��(���u��
���}d�!�~����o}�l_Txՠ's4nA�-�y�B�!���ј��f[�wcY��;��!�=�������߰tF���4*����ȹ����RG����J�b����{�����"�g���-ο�K����Cވ@�k�O@y^"2�\Y�'����P���NZ��G�'�xW����9�m[�8ee����V���e��-W�u!�-h!(GoP��;L���K$g�i7�����X,�qZ���a�*9��ư�'#�[+����z�i7sW)Xt���
������4�9.\n]S�6�LJorQ�������d��H\C������kG
���n<W$��*��aDH�j�6;�y�%e�bnX���W-7OA�H�5��xSH*�Uw6ߘ�e(s����b�(k$R�����T7��6�� n�wLxI,�&IS��$�uOS+��+�OB�B
���pٻ�zf'v_|���������7_�j��-O��9&�)���_=��uU��'�����E�u��ξ�ӝ'��h�����ny��n��O�������1K���M�g~����o}�Y�uO�4ӝ��%���6�>M�����2�q�o�Q����!�T��1����{�3�I~&����7�o�G�lyfᏆ�\��\�9��eÅtK2T�2Qg�C
���[�V�ԯ�So���pb,���Ν���cJJ�]Z~R���x�ya�څU��N��v�JS�]�uO v��zz�q-��!�|���Cʛ����z:誙��� �s��<g'��Uz�99",$,,�r��G{�EKܹw�J��������Ҿ��P����n�җl�qH�e�(�d����&'[?�ȭ��b��o�H�g&z�uO���Ι��g��ς�����ձ�x� �bt�p쌱 �0���R��Je��ny^z�M]d��L�v�\+�pc������·d�V�ư��/��\��P8��ͷܰ��j����kW��{;��Dc���&�N��G�n��אR�գ{��c.ճ#Ka��Y �pcSccmy���}i��W�������_ˡ&��,��Ͼ/?�^�ۻ��Y_WQ�����%mR��xzy�Bn���ƩR����[>�W	қ/�C�d>��&!*\�4�~+z�����=���,��¨��Vj�E `׋Fur���íI����Q��[.���Ŀ�F����
�/^�ۓ�����I�����Fz|:��V���Ahu�~f��jؠ�.����%y尃�`]�m����7{{{Ӛ��WW�\iܟ��B�[�\h��uxr�)3I�I/sT>�q��k������w�.7:��!B�Ĩ���뚁2ܥ4��Q���|�_����Է꧸�|T�����ol�g�]��n]+���[O����� ����'�f�D��e�8~�>_��X]_WK����<*		W?z5:?̫�|�����[���z�n|��y�+�v�XL��oX��?��;���?�.x�K�j����e�U8�o,���a��}/�v�uV��eDe���X���k��!!�O�B��C��@JJJ��pyh/\7����H�������A����A+�痢������C	��S��W�0I�e7�GG�=;V�����C?�sZ�#̩>Zz�~�2����_��f�aׯ_/{{��#�PF���W�X�3��ʒrN�p�?^o�S��`��,�y�h����C^
�Ğ��^�t����L��.�ML�9��
Րh��o���$�ފ��!ϕ�&�Q�b��郩6_o_3R�q��rrr7�a�$!<�UlM�o|������:y4����Н&-u��3}S�����i�)Qk1f�����D_w�o&�?%��䱀�tD��q�WS�3�:�*_�����l;��y��L�; ����/ZE>��~f�q�~�08��!w���cv*���'��?n�=�>�c�G�����KT�o��Ya��Wѹv�����~x|�Pa^;�bn����D���ˏ^R���߰g+_[�pHg���S�Ù���a&�W!�:�t���C�߲[�a�4��S�<:�~�{V=u,�Q����1��/RW~+�o8b�y�S>Ҹn���Эg�*߯F��O���u9��A����~��H���//�g����������h[�l�8d����-��&�� ��CT��U�m����0颇V|+�P�
"� ���Ϳ��1��}$߳دw�a���2�Ҧ�	��>����-5��������?X։8���AHI\\<�a������|e�L�'fG�@����ս�Z��(��t�%�o{��B���2x�?�A�Ws�B
;�_2W���2JZ�j�[N�#�y0j:��+
�}7Xd
�ѐ;dA��Sm��	A��/쬕ƶ]�;z��O�o�ΐS}�T��vߕ�/)>>��ǯ�3Y�)�E��WU,���oS�bj{�z%5��9��rv��B����'�I;����Q��.��g��W��x��V6����kO�M���U����.�A��c�AH�`;s?5� ��Ư�g�~��e��#-8����d��d��iB��曁H�R�y��zR�	2��b�cg�[��\�yV�[����Z~|�mh�T�����>X7���`�@�]h1���{J!^���]삽�	Y#��4�ؑ?� ##����>h���v��|Bcӧ�S[�W����:::N]��[g���p���e���`^�����`��oblO�̃$����c_M���uH=�8s�D
H����M�<l'eNZ0˺ugt��(���U��-����l�01�$&|^V��K�f!p�1��*baL��ofa!���ک�6���F�jO���S(���TWRRʙ��y�_FR���pj��TFKe���w�`Q�!7;���<&��j�e�~PT�3;fϜ���b���7�AT�:�z�-�:�¦��e��lu�8WC�WS�+�ڹS��׆�d�gޠ��
�b����}�1����M<d&����B�02F��r1����b����׫aEO�GE�H[�D�����X��Weii��� <����!���5��zB�3L��G?�,�8+uk[uƔwW'/d��f��U6��5Բ�����M��<���m ���@�m`��������:�	�=Ps�ꔢON�ѱ�M�Lm/p��Eu���~C�ͳ�����4׺C�-���mG狫l��e��O��՞��v��[@@�3V<��"n|n��7��^5�Ow��^��T��W;<k&}�#���Z
��b�Sk�ng��&���ޡ�Z�f�=��LU�6��DA@@ +�a�d�����>���"XJtaI:M��[.���l�����;�� "Ce�A�Ҿ�QYBIXUU���Nb��[�	:T�Z����HTD����Xw:��^��K��rrvF^.�^�k���o�����69Y&P�l�b�@u�Z�f���a�ϔۚ�����%å~3.	�o��~ۮ�tmAȵ�C�,$��͠T�*��׹9'��#Ve��aA�����0J}GubcD�r��B]���{����Q�"'z�N�n�5�F>3nߕ���YWj�z���y��<� L��qC�9��.�ª$���Q�o�Ɂ�W���'��{�P�Ҋ�N���e�[!�޲Nd��_�[�`/�33(���7/
;�xm|��d.<���;����^�ߍ���e����Q�pAx�̃%���X�	y�_�p*ڭ���-;�S2;P��ǉ鰛��-����s�6mS�+n�0�J�Il�<�E<Li��+��i ����C���e7\��0j"�ςx���-��)������|�:�#�|�u��;W%��b�.7Zo��'�������q��L��FE��m)�z�s&ff��kF��~���L�8��!��E���Wj���q��5{��	t~P���KT9����ּ�� ���w�3Ce�l�KC��j�z�m�w�Ϳ�1d��E��x��c��@n
X�S����K�
N�M�B��[X��[������
���/���b>����s]ه�������[ϴ�#���q���[����a�*�gvv��j	���H�.�\23���Ĺ�T,���pو�xi,ѨN.�%L�[������:[��8|�����6���Ph�Q��Z������>���Ŭ:�H�z�Xg�u8��چ1KD��,%��
��1�g�+�φ�w��jJ��q~������x���W�^��[�4pD�'�~<5M��+�&"��k�T����XZ�EU"RZ~�|a�S�]d.�َ��^%���c�K�DR��/\F���d���+=����ٟ����z%��tؠ$:1'�9���w���.���d'�+��,��F���l�����gx}q�a�i5�����	03�c���,����u#j?�|�%g:q.�8��C�xؙ~����$��z�y�m�ۉd����)G%"��~�{�f�ʵW��?��vd( ��M���ԅ�(�{�T�1<��\q�yE�%�ڿC�N����c+:W��*XPD� ��o}3�}����;��i��`����N4��7|�鏈���Z[[_D���$�NZJ�$T���l�q�������h�T+ՂB�X��d��d�ر?���aԞ�[��S��0m��K�c������H��))+�]s4��'Q7��ܹC���j�>��IG�ٯ����L� ���lCC.�Ҫ�;K��V���
ſ^�J��繯�`�o��@�;���b�g�<ɻ$vL�����/���^UV�'$%�!�GJJy5�A�s�<�m�mN_��u�Pe/N^�%zطׇ��q�^}�j]���W��u��ñs����}`{AEG� �<kc;Z@�ƽ�70<��Ǌ!���K*q�"��ƴ"�A�o^���q:�wtR;���OX�$,`���v!�U?�i�?Ry#M���rxV��%dI���g��9W�� �򿫖#H���c�}Q�.]�'��3�o/Gi��o;[{��a�w�������CۻB�������D�H�*Jض-�JrՖ"���*rfmɖ"9%��1*�!g#�$�!!�qr�a0�1��9�M����y���cwͼ���������u�o���?��{Fq�۲�6ɐ[����Q͆���_��w2l�t��U�����wp�`�uP�}�;��"�U����'�7�e�l��$��reưn�S	繤� �Dv$v�ҲIl���j��V��[�$Iv�I�LͪȰd�Z��|�yk4)�%�&)��&gK�G�T)L��"S�KaR�[P��ZTBB���U�ؠ�����F{��9��n�G}��y�7rݼ�7�q[����%�ۄLR�Z����nuX�9"tL��<��l��?�;SWWw.��л�u����[)�r�'v'\�������aEl�갚'�J�v��O4�c�<R��9z��a�MDD�I���>����|�;[�}�i�!�#��t�)z�/|`w�%�'mk�Z��?�[��u����Pۖ�5�A�_��ohi2�c?���e���T�؞c�Gy����!1���BBB^��wߝ��8��>���^�DT�0�-����ǏH����U8l꛺֊W��P���%bا���MW�u7H'�
���I��	�(x"�a�f��ׄ4S�?�Q��������a1�̝3_Uh�߉H�[� M�ْ�K2}n����@xS�91����OlJ:��K��,cZ|�dE^aQ��c�U:z< S�<�@�G����r�*'A}᷋�{�j����g�U�_�	!�?}ȉ����kV����
�a�� QI�����.#w+�����X�C�wә������VL��Y��ƍ�w�U�
��)ҷP�vO
��I��G�?��ץ�]�D��M�h�_��D�qk�n1Κ�(!�"��ޓ������u��om9�X�G��,5gΣӳ��dI�� 
G�Ҝ��֖�껆�R�� �>�a���`?x�r�.���~�4�Ϋe���5q��ʼ����Àď�~' }}T�:~�鹿��7:O����p�,WX�����Ŧ�n�嬨���|,[�dx�fw�]�7k���p���v�G-�MbE��u"9i�{��?��]Qս��P:�e��q�*($���-�r+ч��I�
Õ�����Kq*�n��E��q��m�{Q�w�yU�ӵ�۲z<�w�x���*HM��@���&��jP�k�w�� �X��Ks(��}��5���jH./���R��������RRU�wp|�(O�gn ��tM���������_yZ�*C�d>3����(w���;�|@��)��D��~Ke	2� �E֟#wd����+@��)��ΘxQ�2��Xp����k�ь6��~"|N�+i���fR�5�e��S������"���i�퇔U�!Ł
?Q���"">le�KE�q^Fg�J��}4�P�{缽������Y Ȣ�1�U��Sby7�;����u�w����\�EN��V��_�|� ����U���
��zm��cY&���Kn^���z�֣�¾���7�HOޛ7�������^����\$Z������i&;I�Zf[�������j	m��HYS����s�]������J�g���6��l÷�h}��a�۷Dn�T�����޽��C�f�=��l���9�S���6ӝ8����w����M"Kv61�2n��t�۷o�K&L�2�*w�����<�0�o�a���xY�=?��G����RO��ݻ��ѕ����g�b�؝���R$5�m��qAwܷm�ڿ��0����E1�jv..�Fqx]�Pӆ�ow;��0&'%=�e[���Q�}��������	j�P��i�4��S�f�䫴�3o��xм�Q���}�<'��>� N�o�d+-�(�i�w�%xL����4X�(����L���u	Ijo"ᘌ�KMi��כʫ
��rw���� F;���xk�
)�x������G	8���pf%����NG�:~��Ї��|F��e��1i=C����e�=pB�����,_v���X4Q�^��I^[E�1^
�B`%����v/�����Ȓ����C���se� g�pO/E�-}h�.M�+"{��AG1�1��tl��	��:;�9[��p�֩�P�å�`,;wy�]o�O��r^y��gn�3�IaQ��C����zKк%�t{~4��;?w���,�s*T<$���g�Ǯʱ� hi�?m��\L����i�5�<ĳ�Ƒ�F{q�v�3�W��[I0\�ژ��ɺAV�}�Jٱ[\�	�wZ�����_���� ��j��"s~,B�ЉP��b�
��ݭG�bx�~o�:P�{Ϟ�����[�>�(*)����H3Iy[k!C��9/��ad/l[�0�g^:D�	�p�R��J�.?����D����]��VSc�7Vh�"!�P4�4���\;<�֧�V�&""Y���#�G���-���L��'�vE�4������i،�.��]�/��&Ӎ�U��&T�]�HҚ:^8Q��ڞ{���N�q�����c��T������X�Q�x�pKC��$����7�BH]��ó�h�}>��r��q��;7^..#�X^�(�?����r�͖�/��zс~�"z������UW�Wr���7k��G������eB�]l�~W�&��9��w�y�ޓ�c䮲JjFl�h-!d��m��T �B��������kW�no/�f-:ƂY�����H���5�hP�E/\�ƁO&4�l&"@��!\F5ҋ�>�\�v�P���g�� ��if�b<��^&��f�b!9�I%L����Jz�N��oL$טe�ɀ&���������'�S��G�P:N{���ṃ�=�<i�9M����z$��nJI�.�=}�9:��l�V8
�6C�(䏧p�^
���CE�a�05S�$��e��4!S&L�g�MS��|�z����
_�.�R�bG�>���蹡1�A2�XL�!�ѕ��:��d���W
�2Bh�����[���/��YR�PS:b��K���p�ɇE��#���F�ח#=�¤�4�'�b֑���^3��ߑ��ŚɖC>����׉����c뎚�Pk�T+�k��{B�L��	�8o�sap�����_��5=?)�6���K:�K(���z/=ƭ��D1�W�n��
�J�d�w�?�	3L�3�3��(��
��{N�x<q�X����;����!)]�BJ�۷��p��>��"��ҕ�T`���r5���yL�Ug�"iI�D�)���.tR���C��*�$�=R�?g_2r�?vK��8�t��"�>QRg��^E�����W����U�V9Ġ�R�-{��O^�xaF��{X�F���� {���t������5b��6B+���c2����2��uBd��R�Rl݅7�_��%��H2ZΕ@��b�8��	���7�D�-@�v�ؓz]�(�k�O'�ĩ����Q�k:�f��?7��,��a0�3֊��$l�J-�	��H�[����F3sHx��2��,���r=(�?j�Ry�l������w���9�J�����v�8����l�G�ք�®y�̷���R,�����[�ub����3_ Mr^qe���	�����7*�O����pY!`������kϰ�G&F��T.�p-��m8����c��%�u��[�m�ǚ�1��%l�����X��!(��)�5z�DxL�m���Bn�[ ������{�p . Ћ�x�&��$ڪ��Bڴ�3ӳ��=yD���g��A�<ܵ���ܹ���Ё�{@j��$�$�`mq�G'�FCѧkJ>���K�����%�O�0v�^P=�mi���Y����F%2	�DEݝW������A���tc��������
�;`�\ב϶�O�4���TmQ �=���NJ�Ƕf/I���rS�K�������Y*Ɉ����9�v�F�1���íq��;4�?T�a	z񬴤��&�1�N��O6b����Uz�~Rv��U
��|5I1[�%���2��HҚ���Lmξd1.�����]M�:�/\��ز'A>;�g����hf6��F��9�@�@�+��Qa��nKDE�뒁�������x��Ww����RR�8vT���j�>�Yl�e����c�o2.,�����n�`9�m���=�[`�A���Gd���ź�1�)��ӧ?��J�e����ŀ$z�Y�<�2���=�������&xwx�A<�4�����`��8`	ߒ�g��ooRr��l��o6`DZ�+�G�-X���a��c�wUjhakJUR����VM0A֏�}�)CM�@�Pߐ���J��q�@q���N!�M��?�f
"�ղH:�C���U�s�g5G�E�� ����)�iY*���Y����#��u	��W!��c򱱱������чӑܞ�	�����0Y��H�{���=������:�4�"�e�J�u�6��$r�H{�\uw�4������yX���7��?�\�g�k4O_[���=�F����_)ϝ��Ґ8�J��,˓�>�=^�84����K�����K���}ߗ�}��%���bߡW��!����c��|x����7��Ƀ�<1��5	-%�dڵD%�tx^�4t]�i��abn�-��R7_�e��Q�.'�ܔ-6� r�蕑	2�-��Z<#�Z.|E��z&o~B����'f0��.���+����_�R5�鴾KYWd{b��T<8O�Έ�����uaz/4�L�VD�V���Ҩ�r�{��{�YsI���o����}��K&�q�2�Z�D�4�D�ԕ��~�"�~m��2r���-�A����EwO~+g�X�뻥%��jJ�v%�?���8��wxP�~��[�#v�c+8A\�8��a���kJ�Yz��U�%_��+qb�`WG�W��jjN�eq����c`���������Q	�aJ&�t�(RJ��&���ډ��Z߆�,�s,��h"�A��d��ݿ�-�d��{�-W��M7��$�q������sW�Ab]X�2��1�.��O��;~9��h���y��x5�y��e�ņ�������?�k�@�ff�J*��dPC�Tʗ��o)x��R��B�U�p����:��?����υɅ�m.&Ο��Y���@��q��R�"7�c�ȩ����ړ���b
H�^�xU1@�ZG\}|��峮���^r<�5��^W���F��m+6���Y�q���P"Y���c�ڨܳ��E�t�E�g���1�g�����m�� �^k��E����9�}8?��^�n��s2�� D�A)l4NWm��qB��U��>��Ay�_?��s�=P���=�G|�h*���b��&�3�a 朗������c��l~J�����u�n#Q��ܶPo��3�U� {�#�Gȴ�?P[	�^V�St~v^��\���ʡ5�;�� k��f���?������Cb!��b�� �^WAI��-��"Y��Ũ�4���]CͶjT`��q<u<�˅Y��H��F��d��+X
�����4�c�m%~JG���#���T_��R���c��*������)�OcFZs�[ �&��:ۖ��goJ8*`�\ŷ��������T�l�x�
!n�/Y�5'�5�̕�5�3I�ݯ�*)�.X�nuZ3ڒ)5��������� a���0q�n���Ua#�&ɞ��'q|<�����۬��x�l�p���iX�2���;xv�O�j#���I�����ՙ��:�j��N��bC�{gL�VJzO��*^}�:��i���c�l��Ov"~��٦�7�!$?zb��}��Nq�p�5��h�q�k���Ua��P�+���h&�B�Tz����<Y�u����V��$�����))����j8e���Z|��(I��Rs〙����64�u�Om>$0|h�p����3�
���M�SٽxJ�+�߉q��!�g�Ծ�_F��yn ��y������;eee~�����p�A���3���CTJ�|��*�iaD�����53�Ka{��}|��N��������Rm?t����]��aX)b�7�J[�CBI��.��т�y�"����R|K���&ov*bԎ�7�J7s��X�l�Ʀ?�+�8&�^�暩��3���9�3�XS8�:�A�t�_��<ZV��H<�|��9�؋Os�F�M���(�%z<�]z\����OU�3�w��83٭����_سj�.�0`i�Q���R�	M
�~�E�&z6E���A�c,p+�@���7E;G,��_
����3���jTz�	6�J@��w��D�W�t�5��yqBV��F�M�%}n���j���{�.��Y�b_��N-��0/«����<�!?k��b�����V6�A'~>��5b��M�.Zv��(�1��G�u��A��eS>_J�>;-�C;���K��}�ơI������ ���k�/��� 
rW��M�/����9�.�\Q��y��5b���'h5E��E��
]c�ln��߅`N�D ��H)4�"N z�K��h��k��u����L����B���lJ�LR�y��>pa^x'W���`'�s��)�� ��z~Ia�ȉ����z������+%��܅Q�c�G���E����
K��d�)�j�R�mq�`��/���-e�,�O�~�z#@�x�@\-("�uǥOπՎh4�͸��Cuk��7��7]h�v~,�U��u'xS��o�ͦ�)�NW��q�k��~ s��c��\(�ьiH::omcl �	�����/��#�6��-�dI�]�6�+�9���5D��1]��dM.j�$�YR��z]���!�h~�����HEn��WW{���͓~/�ۙ7��֐72��E[��EsS�!|���т�ePWL�'���Kth�v�f��>KF$����w^d:X`(c�8U�>w�\���𑕛���=�C�g��)����4}�W�+� <�"?,��� JLW�A�g��P�Ӎo~G�S���z��kE_�]��>@Sx�h������gh6�?�����BZ�&��O�;K|m�V�)Q�#��+� ��%$r�y�s6��P}��W'�C(����N�Q�v.���X=�d�c%~��Z�p�䐀�7��ZLTB�F_6,LV��7�^�m۶��;5:M���I����	|p���)B���M2n����G��]����im�r���ヨQg�ɩ~bi�� �$Q"��ҿ����,8q�����`/��@�$���{����L������^ȤDߡ�����3�ϜUpV�l�3�۽B��{+�l��˶�zQC�����=}�D�<�6��M�"@�X�Ζ|���|��̭�Z_Z�YI��ny��6��O��}&�&�g��=�r�޸�����}�=���ͧ�{j۴�"�j�EרkU�P#EEųZ*�6|�-�����db�po����BTZ_��7*�wwP�F�a�͌���qB�J��� A�A�9(~�a�	u�^W@dLL{OK�PZ��ɷ�	��6��L�niw#h!���2z߂u��Y���	�_Ť�?��̔�F���\zB��P\u��V��E~~�»�a�:�S����.�J!M��/�%��[��q�Ͷ�txGƈ�a�鰲�ւ��K���̯ͮ�n�Y�7�m����w����&�l��z�b741�@�G�h�iB�KX����o+n�V����ޮ�2,���"$zI�8i6��ܪ�3N�c��!LTRP1DR����ޒ)�Â�:�7�_�T��r�D�Xz�@"���eg����W"J�
�p���T�L)�� ��TO	Z����׷�i�>oo���zaa�x��=���'wO1055��`#�����p4b"b�-��q���Pk�z�A}$?��Y$Q�ѭ8ey������	XR�ޥ��4�
�
�e�t��ǿ@����c��t�/�V��ų{�̙�PT`{�ӽGN��u}���ʖ���jm `�Z��x~��Z��	�~�cƗ��m�ջ�6��ew�d��i�[(�8u<�Ȱ�G���9*>�i�����A>�d!�)ێ����>b�[G
 �/���"�Y�0�Ë�>��9�7u����y��9�
G^�5��=$��6������d�Rm{{�x�0YY��IJJ���g[����Z������G�G���iaY�:�#M�5�8�ү�,���0n�ѽcg���$�'-�+$������(j�v}r8O��[�5���A���yD����!zvjdp�B���W�pt?)9�l�K�_�'u��D��MJJ���*L8�^
O	�h���p��1��)��/i�e<���0q>�\�
I��GL��&��MiV����׏�ݻl �l�C�G������7�?D�#U��)L!���"㝮�ڌ��}��124��$�V�wOF�������9s��ɉ	��iUMMM��"S��teñ7��n㚈]xJA<���� _وR���e��"�����N~h�}�K�0�h�s� N�_x�����m�ŪO*k��#?�+ۊ0O�'�"c�g�I��Lo�9K0��}7+�)�J�^JjXR*6@"AtJ�`�啔���������7uʙhJ���{�|UMM�0ߢ�#Z���Bbфր�KiyۼI^�ULr���fR�h�:C�uL��6e$��%�Q�|�$}��s��K9Nc&�����l�Ob����:ȷ�^���҉<��!�����׿�1.n���&oW��tB?>� jW^N~Ri�ԡ����;x�ͅ�*Գ܁�e��^FπȂ��`Ӵ
�d֢bͶ��f�rp��#0FIbN�c+�.I�i�zpP+�ȼjt�h��S5���_��S���Wd*�5�B>�oՊ�V�ytI�$k2�$$$�k��-j=y===�	���X��ӥ%o���ett5NMb��}�4��k@�X�2N6����}��xd�W__�Sw���1���(�� ��aꟇ�~x	9�Y����]^f�$�n�%nJ����~�W�9׈�~����ˇ��&͚=:aO��7�8�jm�X58cK�Ww@����FNv6�餽)*�ΦV��fi<}e�e*�^,�f�Άpۖl����a�]�h��D ��H[;VH�ч����:����5_�ֈS�3_���L���������u5������e��Aڏ:&�Ԋ:#[W)����U��5P�g�?`M&L�7)�bia�K�w_��d���kOL�|!���x{���0���X���>d������=e1Q�~�ʭq�� <ݣ7X��75NQ��ۉ{N���`_�HhD�!�:4���UX1�O�&)]4�<*UG�q�C�������l���jf� =�B{5�%:�P����S��E�{�P�,IP�蚕;(S����a�������<��}T	��K��Q��wUe���%:;Y<&�uCݾʌ�?�)���ʣ�:���"���B��G�8���$ }�W��*$��P�H`*oٛh�eԩc~�%��������-�11�uιD,�'��Ib@��;�]fGr�W)^��w1iA��('0�$�aZ����L�j�,ics����O$�Q+n�tttdyPοjY��?��hm�S�}�E S�B�	팄���ᆪwq�1$���x.��s0V�A�b�{�3��s	��3����k&1B���
]�q�*H@@L��(~�A{�6��~��g���A��Z�K�z��*�:(o���;�=�Q��'�1Z 0��\�*�O�r=˰,��#�w�5Y\\L���������{�3C�Ve7 8TB���dz.��˼�����|Q�8�9=�.��6tL�e]jJ���e�A/�F�4y��Ը�H�w�NtP�݊;���u��~��`z]=G��%�\�9�nˠ��W�OL]{�mj/=Y{2e�c�z��J a�hS"�	yyyYׇ>����8���%N�w̕���!�!*�q����; %�4#��gϦX��Ą\��(.>�e���g��۫2Ԁ�/r"��ޚа��'�t��H��w�k�Y9W��JӇ�� �$��S(�`q+Nfbۘ��	BHGi�3�ц*��2���S}��2�ɇx��=Bt�L�24��ZG�)�w
Mh^C��:���Y:�T|1�������^ՏS
����QTTt��^���,nˇD�X>���̉�Ë|��<�Cx����[b�+ѷ=F����|�C�f��M()s��������_�����^Oק�h���������o�<_X�K>�Q��B
*�s����$�W���-�Y��^���AF۶ ~�]���v�m���Z��4���h����J�b2|�U�g�G��߅V���� )�eT)�K�J���JY!�K��W}!�:=���xk����؋�����g�h4w�6;��_���08*��𝄂�b����8q�k��t�yZ^�������*E#���u���G�ſ�S��cw�{@�!%p��Me�V����ȕ�ō�j������L%,�,���ic[&�����Ar��W2�/���M�2�)%E��H_��LO!\�8�I0>A�a|�T��AUc b���{Q�&���:j���'{�o���zʣ�k4Oj�^q�d�D�A�1���U�i�µ���Y�����z(+(�}1��jN=w� )r���	�QX�~�1��t
f=��U����(_��R��o�B�:�kܒ �c��(�D�u)����s����~��p�M����<���?J�v8H��1t�\G�"]���k��m��B���W'���O�����4_��S��k��^��k���H��z�[da��7Z�ypt��ԑ̹_,2�C��u���ȓ�*^;��mԁ��g�<�!t#ȾB	��1�'��o�N:�l���H���$�=O,e�R�{��J�`h����Wd��8Z�0ɨ�_]=G���f�����bz�\[��8�\��B��L8U:�	��~κhJ��ES����L搎�K��ˑ0�]�R�G�V<�Ӳ��x9�>��\�o��Ё0]��Y�oI��447?|pt�c���p��O2�E��������=x�BP�����y��>������e c]&��F�s�(����l�Ǐ�qG���FVn��Ң�M�q�JJ���p���ss�j
ݿN���tL ��}����M_���=<eN�W�-u�����l٢�/�&(�D���ܿ�Xn�� �6G-���+�(�p�֭�s'��4��M#���7 gAj�������q�Tr�dl�����Qjr�>���X/,h��'��^�s���������x�qh2@U�@������3������R;[xޜo�-u�Ѭ#+�~3OQ
����L&�"=[H}��0:���n1q�27�N��:��Бq{c���K2�n}�g��#^�H���{��ѩ0�wttү_L�eY����������7Dn��%�}Pe������'-R��5���*Vg7�)Z~u�F����Z>s���<�g��Fs�`0��6�\�2��D��s}c���ᶈ;������=�������]tӦgo�rr�:
�Q�wϯ�^{N����{�>�m����[\�m[ο/�r�����S�㚋�.��X))��O��H؏������1=���K��_1��֬��_�Fxy�ԟ`z������8d�Ф����Wh���b{��Ǐ�4�N5:aQ���@���[�Ň�S����K�
�����/�9���GY~y��A�n�v��ԍ#\�9SW_p����b�J�*�h[m��ۊ*v�!�}�rɔ����7Z��z��+�T�	qzt@dn6
���:tI*>�ky������]]7j<I����!{�X�^���y�B�mw��`�J7�7�w,����QLL��ղ�J�?:/����i�� N�2� �a��l��k��qmڞ_W��]��F2�8���Z�j�1��#�>%H��
0�_�X��U!���û��?��7{_rV?"�(�ʾ�[�U8�ejmw屲��8���c�G۝��Ŕ�&Y&9�A���g��"
��Ų[��xL���r�K'�IORrrC�A��U��O`��4��{���S��T,����D热��wF�~�+��U�na}<=Gv6%d�:�|� ��c���PÃ���U�a�D�u����x��������<��(0�̝Ma7e��;�v�O��z�hO�6p/�~�~�sX�d����C$���+q%91с�#�<�c33���8Y�X���'���t(�������qR�4e3�8�ž�ax�C�xC�0V�?;\�A*dji*)u�Y|���K���R����b_T��'�]=�I_f��ˈe���O,�q|�}�~2�8�}�h�V9N�E��M]�q��/�3]Ր��j������e�wN�c{��Gc�93�n"YUfp��Ņ���uu����h��9�.�/�{�F8:0�x��av*�����-Y��9�A����9���J�*dA�.���
��e���-ޝo~�Z>|����G�d1�B��$�-Zay=�)���-T�Պ�l�\�����]7�/AV�֧�E]��j�9===��ֱ1GzT�|NfF��)`!����B6��0���{��1��(���gk5a=�=��V�̻�f��%>$2K�C�,�1E������^\f�x�`��-A����y,�?�~$6����Lff����3���$������c`d$��Q݋�h��644�l��*�u���W��7v��m˯"�ǹ���@V�o�=��
�g����)$� ������h��c��5bx�G����VX ֜{��e1jZ;L
�����_������ֆ�$#��V:�]J�q����<=���J2>~4�24�
���F��p㽃4C�)��S�ZQ���u`N��X�Fv�gL���[f�W��q�/��q7�?�68MM&^��CN��?*�RR�2���SUF���G?}z��	x[��Z�>�^//�/$�Q�;���=!�/��'���)Ŋ���6�Ħ�L�j��S ���_k�s9�c��������>u�sKɴ&�u��W�_�)����>��ĳ,�b��B�����%����~�|�A�y{m��K�����%���l���h޿/�CY1эe�7r����ݢu��(�j�Jإ��6����Q s:B�Ӹ��0�>6�\���Ã)�^�Ț�s���U�q�����,r��|��w?ȧ� ����އΧGY��y7⃴��xO��@���^��Npbb"�����k�X��<QjN���좾�{��!��٪źH��P>t��#��<�u�X<Cb�s�U����y�2�Ռ+#�'�\=��Ѯe���'#�+Z��&~uO���׃�XLZ���%�ƬZg��,�NN����:��kl�-��!��7547����ulI��)��X��p[�E���k��t�"툑���n�'r7j|������$QIDg�;D��_����Y���Ɩ����O�ho�%���:{� �0 ���=ɕ�
T��
3����f#������wU��{��+X9i�]~nQ>�ȿ>�8>�����8�Q���5���ʳzgӦ	�����坎~�3��Pddd���g��F�U�@���/6ë;���X$�~X���bq8L�fGى��5eV�x�����I���3�(8�y�KUF�&'6�`�ݮ�$4��'�c/�jC������D�3��>�l��M��Ɓ��C��h�=B~Y.��R٤ͪ&��E���
O��C�\P��ei�� U����I �k�h�	(��#�I��O�����Z�����{`��'.x�n�99������3l��SK��ㄬҹ�b���SˊP�5�Jxz/ Y����σ��G�|��A[(������Y�Ȳ|�\u޲��{>g���N1����G(��)�%��jbD�m�E2ca�|���vb�*B�����J�U���7vH-��M�������YV�D������!���uj;>rⓂ�;@�� ���a|s`���B:��|��]O�oow�f�p'�n��sZ����qM&q B�kE�N�c�|�w���޸���SV�A��΀2�9x �ީ���kE��).��\�ѹ.x�D��g'B>���c�+1��`Sw �:=���e�'ۘ5��9�+}RBL��0%���@US��r��v�M��j̘d�[���0=R�J��?)E��!���g3��y��G�j�j�{������Z	lb^�b�*v��m�q���|e�C��@�h���ȥ햇t�AZ�/�xw9|e)1%Yw�f

S���U�۵��Y�rn�4����'N�/rO���ư�"����G^�+ͧ�y��_���ZE�N�����l�rmKK��s����������ڎmd�OnͿ�����Zg� [qkr�c�#f�MrWݰ���ۚʌ��"������ZP�w������+�����.�6dr2���S�Ɍ�\3�ڭ|��$�-Z�qң;y�E"��e�r�Wh2e���,pu��a[u!t*�V�0�x�J:�}�M��y3~�-�H&	����n`OW��F$�8ݴcT��["��ď��Z4���I�OD��$�jj$��t`a.+�pqqI��,Y��֍�ci�E�=��c��Ȁ6x�;q} h>^P5��fԝ;w2��R�0�cg/�p��4���ɬ3�3�L1D��E!���j�[�Uxג�6a9�Qt��B�������,�Au�	D�~��R��V�>���wf	�HqO�\i��Ջ�� #�����]�;��KMM����HvH�����6 �Y؝����uuIw;�.���]��g�����$��x��u�]R�X#����������Cw����ܙ��Q[�.�����w�b.��ʎ���&�������-��]\�<������X�PU�ӧC��W�/2�#_KL�XS�ڵ7��دs�51���)w�}z[�f��}��B1W�}"�i�в,x�	C��ެuqI�q��(g������!�@���$�����f�W��}V�|A�]�/�Mp �e�5�M�
R�-3�������D���_�X���F=|�&V-"<Ij�G$�Ś�� `�u�OM����C�\�Y��9 �����Q�-:Ʒ
/�d�M΃��sH�B��2T?�ᙠ�@�_t��3�wff�����3z}	��\x� ̍�uw29C����V�#�ԍ,y��	,ec4�M��������sr���'� ��h�ʠ&�۬��3����'ZW�Q{�����Yhj����C=���j��5��B� ưO��8�ԥ�Ԣ�������L�EA�ߵC��.|��g�T�����z�(|��ia�q�'ZxJXo΢�l85�����4X�Vja��K����P'>��T���
���H�N,����|��ߛ|���֮��t6ts\MZm�v*ޡMVa-���K�
2u������a��z�0���{Y����5��G��5L�:����HY����ҭc0��V)����4`��=���;���������eNH�S�%�<Q�
Qa��<�[�����kd��ׂ]�c1��r�Ζ2�xI[�T��ĭ�X�q�9w�F��z�KJ�E_e����}�Pe�g�A/��Q�:�mvxor������ �ξF�ˣ��J�G׆;}�ӑ3U
���'VK��w��D�����T>��{��E7�@���ތ\b!t�L��!,<�@r]��!��wG���/S�"P�]Q&�Ti���x��B�������0�2�H�U� �ّ�^��Z�5g�F?��d���-���utuu�0h=���������_nL$�5���ųrr�፟]D/HWW-B���)))䌃�N
��)%99y-u�i\h�s�<���;��n������>\uɐ�����^^�`��tE�M���tkvI%��f� ��z� =o�=YhO�7��WI%R0��K
%���0s~dL���pYU�j�@�U��Zv��޽+-c~$�a�o���6,��L;���|�Q���b����NJm�S��5Ѻ""Чr��+Kz嬃GO����Q�"��pНl��`ݡ��༝]�N�5���m۝/����BM���J�-Kh�\pZóg�v�y~kLr<R��{�}/�-���,����E-)�y���G;/�H�����t�����x�`�\K�6"
/$�T�٥��������]�Wai%��[y}36�ː�A�W^��~5�sW;OîlΑ)��"�"<��RwA����^[�������o��ݸ���QS���9	�k�.<�������_g����5n��<���z�T͠�'8n�b+H�4������q�-rx�ڷc�5w!���f������XiK��u�e� -?�
_I�rP�����kה���#	lAQ��!]݊TM���͂�ܹ���%��^]��~���-U�ß�wI:��|����"�Ё����]C��#H�I9W	w����.�/�E��.�4H�Į���#8鸶pҡ�D!pƫA�9^/�?ۡ�d��+��| 3�TR�)}��F;�"��~��|�^���d��|�	>�(oV��:���E�e�d�s���'�++����/��[G�!��LI�#��C�$��Pj�	�i���z�glb3U��S�� +� e�87E�2�n��kR�Hk���AV��vj��v8q2b����.��ـ��GH@�&�nQazԚ��A�qgs�8y��"�Q~�[�vM����o�+��Ue+.N��/���'9��}ܘ-�Nk���'E���������C:���Ч���=��!&ohUf�+H�7�︫�X�J/L��k�.� �)�0�H9Sg�B����o���2�Z̉�f.9�3�J���k�R}]�����]���{"�F���F���''k��;�M\\|0�'p��ѯ^ݍ��Ce)�Yғ����ۯ��.�좸��a`p�0H�wv�;˶g�a��P�]�,9���TFS��}`�"��~;�VQ\�R��t?�rLxĘ/a�Gу��V���҈�5! �I[�4��&����2���Տ\��,na�`jAa��T�n��fs�\�c}A�u�W�݀���D��N~�O�0�5��3+L��񄈩%=��[�d���2�7X7�M@ �P� �S_n�ݱ�[��=>s�����\��o�����Fq�c�)�8�K@��28(3�Uh���+	y}�g��������u'½w�i����N�ӽo�{�R���JjL���~��G߅����j'������,ԒwXǆ�$�ɏ��,���(X|Kr�v�B�Zr2'�TVVF&Y�!�w,��	|��u)����>}��:�0��餫���o��x����$r$$������V��J���nd;]ɘ�=�X,���bi��ne�֓M��?��S'^�����~��T�u��=뇮L��&�q)%�NEIiC~ёn��z������/��~���Aa��8Y�N��=w�y5��alUTU?b����Q��&\�'�4�#���)邥���cx��*\瞔�2s$��z��:�O�Z	���,O��[�����Kp�2��v	���	�OG��ѯ.��Q�SM0�(�~;k[[��II����8�|���T�mvn�j�qV���i�!H!ru�Tc��g�f&���GF9`��T�=+P�d���!��3�F�J��փ�+��W�eݭ?{ɦ=��ű�r��ջ���kz�{������l>$H��gE�J��*�86��z�$l]p�	 �p���zҵ# ����)�O���B?�,�>������bfd���_���|�eB��O��ΰ��\m�Bb\/��g�Ȅ�����m�����'B�6m7�A��|�hc����8
"Э��;H?�D�[P\��(e���ulN���#����0w�u��p�j��eo|]����P	�3�ED�m�T2ma�yq�Zc]�e5�&���������<dTਇ@g�<<�<�~��u�`*ܰԵ����*/�������(P4GW<��'��:��+���aS��@��5��8�G����/�q�(d�!��I��ۻ�%����΍��?&sł66��r8�����>F�@��"æ�o�����P�8Zja�>U�1�Ֆ�xM�7?Z�K�7k������~9�K��k=v�"a���4��%}��M$N��6�>';�����$~��ڤ^���@{���2
55�P�Ů5P��Ne[<�Y@RŞ�y�3@"�уn�5~kBC�̶ZilUHdN�[*�b���+EЬ��3��L@�BՇ�j?�ٝզ��5�(U���O-��R�g��ؔ���D,l��3�����w �
S����y���C����9fެ��9�,�]��s}����;_s�
�(88��]ƹ��2F���q����W��^6��hg׶j�s(`}"39Y�z����,>�ܺ��S���>'�_U��������]ߠ����,��+,]�=��d�f�v�~{\��Q�G���gS���r	����8�@����\�l��a�/l��b��mZy��/&��$τ�	3?Mw�M2��j�^�2z�=�#��֯ Bӗ�Ј�mOXf�7��[�
=\��#ny���nt3�X-���4�R��_�u�{�D�dT�>��2�� 'r��˫��:�lAga1[�f��qh���=28ѩ��(2_�04���&F���;i>S~�z�w{�Y�G\�V��j(�z������+|K��f��r~B��� ë`�JK\��A��%\]D��=z]s]n�����G����s΂}�t���ѭ�֘
��-v�\�
C�s'��A�ޙ�����r��DT"�Y����AB�'Ug�o�&?f��>-E$HS�j×���lAWפcO�A6�8��o>�����e?ǵP��pP���^S�����ؓF��..f�L�IK�r�Tx�]Q��������*��8�h�F3�5�NA>y딬���v���O+�u?��%I�F�G��C�1���僷,�d�kjnE�����Sm>W��L�R��R�ʌ���\����Î�8��&>/���b�ѕ�?���������n�c_{+?�iT�HX@��cȽ�l�?��}]S�2�>lpp����zMؖ��̅�R�7zvRd�����ѻ�������L�8Y��y�������Jm]]������S���N�����g�6B���(��x����۝{�BtS�B;%�=ci/
�Ȯ�}	3�i���Q�+	Y"�u�$ĴX�e��:c��;��0g��=>���s�y�����Z�9)y��q�ah�"�=��kۻ�W>·�����|�����h�_��s��X��o�>ZbseK/���'<˾���g�)V޳���-u�d����)����Ae�@�m/�:�����O^��xJB�E��α��rѹ���s��G3O������yc�Ld+�����/�T��Y|���s���O�J[���}r��Zd֯w��A]��Ш�;L�
�ON6?�6}��9�qf%vvMڑ�lG�9�gA�r�Ĩ�`�zj_�o�_ۉL�����+ަ*,@Lч���.��;�Q��?�`��O��SE�o�������8 D%|o���?s�;t;:ڹ"c`�6<`�b�zz?f��Y�~Q�]�?��~}��§oC����#<�]�R�;1*NV�N5i���v=�׻�v��p�`+�m��sI���u/����[���)&~6B'����:> {(*+���� oqs�}���&h]qv���2����_����@���={µ�0�1���* �ٕP�ʘ���MN 0��*��� �1���ȳ>P�hNL�'�:�Y�{�MPl��0��j�\�d������b���@���Mف1�)� ʷ�Q^�(	.]��#o���|��8?�����$V��e�"_y2�'��Z���)3�w�j�f� ZL�Zm�c2Rv�?~��L�a�s�;,W9Q^\�����Y����J��c����W����T�oG�I'��9�]_<e���jO���پ�dp�_���4��H��C� ,&|�{�3P���F��"1���qt�m�$���BI�!�+��������s���"H����h���}�~���lz������Zw.ƃ�4�	<e����&�ڲ���I��.Y-?��`���QŁ�a�H.�(.@t8G3@"#
������ļ<u����&�.�d�����{}Z� �Ji��R���Ա!@�ߡC�����Mw���\�����^vtw.��Ƙ�fi9�%ր+�81�|MM���u��о��흎4�.�G��m9���xL��X���*����*���z���w>���U�8	�ߏ-=L���-���l~��g�����b����2��P_u��S8f�`�:����D8��6�w[�������
%-�����^����=7"� ����s˱t�����O� �?>�S
p��ȗ/_ZYYm�v,S_��5t�Q���w��b�������Vs�2l^�j�J���)���/f7ܠ��y�ii8�%QB$MA5���S��Ɗ�.�����F+H{�)E��E�r�:k:;�{�*lg{�Y�?/om�D��q}�����`��������)T� �s���3U�ܵ��&�����γU�m}*�U������n=���'Zn�3o���y}��#��Q���}�鸪V)�H����MʷVY�pIe_�}��:B1�Mď��C{&*�����j�����{����A�{���+t|v��im�Җ�~+MF�x�̠�^����P��u�����y�*ڸ�"o�]��DKe�'x����	ғ���,���{9����9�ޅ���_�"�[�t��*�Ш�q���ړW���1qs>=�73��%��v�����	V�/*��/�S��S�=��xq�*>UY~׮A���>��>7�����ub����"�@�Mr	�sg�o��V�q���[V{]&�2��k%���bmL��;`�[�VT�飙rK��,)/��q~�m�ĲD�F���DT��=��p����V�T��N�m�HA"���U��G�m@��e駵Z;��?���� ���8x��(S����q��e�DR��а�dIII�L=�Vl�b_#�6�J�<e�)EZ�[�3��V� j0?�I�Z!M\U�x5��1̑�z��8@&i����^%�bn���Ԝlv�H9��r��}�ZHS��Ю��v�Z"��|�o�붢�Bl��ϟK1���7$��!�d3K�j�_G%^�\?X��x�VUFH� 5�+Hy�->��������1�}��/�VX��rrrۼ���VV����)�lW����h@c��8"��Ex���S]+�?/��,��QT�[Ǽ����"M�����Si�g���M\=�[5D�6~�Z[��d[kW�7�3��x��؊f��/Ű����B23㋌{�F`gBN�QX�����WкC�u��=��ȸ��kV�B��I͑�]�����j�b�F,�I�b�(qM_oAI���o<r^R4��1�r���^F���=���X`�������J��31Bg��	p�M�����1~��t:��X)���x�e`-��o@>���e�?�p��<j��#hY>�o&$�n��s<���ZIZ�K=z�%�n�9$�S�$��V&d%��r~�`as������gff�'�%''�tN�@A��o���Q��������2{4�YI4XUE�\�̼�@@���IvI_/���1`g��z�?����AZ��4[������|���q��X���=��Ā_�V���.!�����?9�����E)q��<�
�4 ��U��g#f�{�~O���JZa[���{�,���#�,�qV�#>�oi�ܲ瓑���#(�lcƑ�"�jo@ ����ϟ8��"6Bru�{��jy�aCd�\��t<U]��q�q�L���ǐ��J����E�~ق�Ns$�yk����'�!7@ߵ��	R�i����ֲLg�'�Mbf����X����nt4�` �4? ~WK!�Y�˗(w��|�k�Ơ�k������O������Y���!�w����DcW���a@���8J�M�Tӏ_=%vV�Zߣ�l�����{�q j/_���V�ٱ� *u�n���������0:ھ_b���?%;�|�Bž��i�޲�Y������oe�@\&�#pG�D���ϾͲ�{zz�`�[	���uM 7_Hk�H�,���!E���@yAh�\�F,ώAo}��1a�I�;�uj�_������<ض�Kϲ��	oΗw u��^�d����Ծv܄Ny�)[�Gk�Ogssdf�V�D*?�E�fV��?P.��W��S;!O䌹������{k	��� �,�m�ff�5�௾�_K���+]�n륎r���oSo����t�̥4X��d�oyE{o�So�}��v�VD���A�Js"�GB���N�������)@�	(�w���Qs��nB�F^��y祝�.��f�rY�\�����?�wD�x�����0�9��JG�3�?2ԑ>}MTT���:R�46�f��ᐏ�^���E����W�����sj���O7N� ݷZ�9�u����K��<���m&2C�6�1i??�◺ku���(Zë���bt���T���:�|��~�Z��`��7�,F>�w'88��r;�b�䕔��g����Vۚ�9������}��u
k�=��@ۻȍ�.1�K*��-p��=U��vR���tn�/y�^�S!��wJD'x8�5�*��u1�#]�ݦR�}��
V��j�q;̨ن4����v�=x]�?<�0!"U�(!!!�Ċ�+��$��e3�?z(���������x(�އ2kH= S�2U����6XvX��-�.�ƍ�ש�W4U�#�j�}���'�:Nꗩ��V���=�������~o*�}��~��/� Ա#-�����d㴭��^jzS��ݺ�Fs�h<���>��˪~q�s�ޘ"�����ײ��O��Ari/��� R��G�Ml|B���ލ�D�L��?���y����d���|�r��
�ʦ�9 �&{(����$Z Δ�b��H��.�=[?2�����h�|���W��Et_ȱ��W&�ox�˝'��Nl.r����O��L��P�;6!y#� Z��X�~���C,�����
9�߃1��Wrb�|\\�7�m�o�?�S>@�_���;���e��Z�{���I-���c�g���j[��9���+Du�
�r�����jOj�̔�鮍����;H#.�Ncϡc╯Al��ؖ�5pSBb}��;*����$��+��K_hx�J��z[���k��\B�{��/����=�Pl�k
�;��9��<F݁�3���c��5���|eE^�"�U)�-�\K2M�����Ɏ��-x� ��>+\���U������/A�ο�yhDwyn&T���qP��(P��-#�
�cmi�_�G�.�gEK�m�Qd
�7����ҾoD�T7c���U�p;���
D�ߘ�Kß������ė����Ϋ�F��gv�:L����e�Y�ooL�]z����(v�^/,��s�ӕ�@�_�5��>*�T��O��ś����g_��N�^�#]yW�䁰ikG�Z�C�7y0�o���}�Smg���pCd�6ψ;n�>j��9 &��rqE�N{���� ���Ț�v��_�]B�<r�+��e���!t��^�;՜T���EH�� H��(� �f��찷a�=og�������a),w�Q�8-������F�_O���G0�7i��:�䤊�
�@�}ܸ����,�B[���= �_I1���jMl#?�feeu�x����ʉT>
`{����@��B�Z��g]��V�5��YR�'�yxx*�sA����/~E�<<��W+�� �2LȔy!�N��5��Qu����2B=�M-�#X��f�2�v����B�~T��i�ǡ�oPe�<䀨����hs�]Ȃ+���?2���5��*��va���w�ƾ,G�M�G���A�j;��Hp1�[E��q���ГrfL��!�@q�L����!MKJ��K�%��oᷭ��L�J�Rir�2�S͐P�*����/_����[ 2^T�5�Y������}�?�i���w3�lY���)���{���t����w�LSzb�����K0��@��d�c��ʈ�ec��m� �,7غ󦙀
��T�af�7P��(uY\m�	�����<	�T�<W�N۫�J�@�0�N���O��f�%� �U�G��1U+��rLBLlǵ�O좙w8�$�|�<���޳i��������:W�������e�R��s���*	Y\~�2����Y��s�
@ް��Sf��#g�f�8�o5_qn⦋q�`=qYF���H�ʢ��(��z��yf��c |�� ��k�Q��bj+B˥� -�lo�� �!���eb4Z��r�)�JP�� ����Vzk�����p��@T"�Q�^��ׄ��Gqy�S����o6�6SDh��\<����i�}�Ė�Br��(�/K-#��`�嚒����������[���1ZL4vK��D-	���0�~܃,��Q�	�1w�V�;@CaU �����骁��Q{��M����sϸ�tŷ���Z���$�E���ZK;:6¢��MI�S��$$���5�xk����8C�yw}qN H-�yiUy#?Θ[Zz.+����.�q�.��>eȈk`'&'y:�~��B���*Pl���.��X��y�\>���O3l�#$+�U�V����d�9v��;�{ڃf73��	T �Uo��97�#Wѐ�Gk)�f��d-+1f.�b1A��(���7 ����h�?	u�!����]#
ߔ�����o�T�#�(`�/k�ǿs��m��
����ǝw�
�7R��ٓ��u�_��$��\�u|�����'e4M����Q.��ׯ��+چ 9������^��Ӧ��1D;��9�NDD�L���۔��>��t�֑���`2vL��~�_����2ޑ6���pM�~��
;���H�
��La�q����U�������X���769Yv��Q�_B� �N��aU��x Y �<F��r��JA�Kd���1̦f��f�Hf��]_D��ja�.�	i��57E�S�|́*b�>I�y(�,�/9�b��Ϩw���Ǖ��[:��}�	��� �Ќre�ra���(+�Arq1�����[�n�o;t�й��h�|��7g���>b�@�-}vo�F���?�Z��J�_�ށ���1\�b��76P:nZz:�Ç9�����s���s�y�SjmåR[��B����4I����Kԟq���{�-�==Pk��1f�_�&��@#�$Qs�c|#}I�e*k�,�.S� ���t�0X�����ED��Y��\��w�e-���)?�R'LK{�Ǟ��������H^Aa5Ԫ�>eòT�����`γ�v�-�e�ccf����a-�N�J�CwA���K�5�봰�����P6ݽ�懃rg��d$�f���j`�rH@�P<=r�f(�$��U$�>��M��;Q���S�ڲ����(ʕ!3�V�qe����9�E���ؾ/qԏ�U�ץ@�$/��2�߁�mvf�g�"f�;<����o��o����t���;C����a͈�OM�s&I�$�yQ��Ei؟����L��)X���v?#�Baf^�s��.��$��@tx�C�pj��������w��˺�mz�Q\�����P��9�(����R\���]�f��IE��'7�� ʞ?��>4~n��G���8��D�E�Y��D�d������;Ǔ���z~���X��2�"���jYgyH�J�w	@r��`�'+��������� ����/3��sr�>�;,.�m�'���/uD?1�r�7�����e�
k�ު�驞΢^��]`��C�*Ĩ�UUU�Ws��v�1~�݌�2���R0Rn}��>Qr6R�	�yU���a���`���uk9h���=���|�yiY��N=}��!�|Y��QR��������_��N��*��w����X�orH�4%�3B�)�P����΁`��d>9иi�����p4:y�N����ϫ�8�Z��766v�
���&�ˡ3<�1�Qv��}���H�Dzs����c�pC8ǐ��T�� ����f�Ƴ3�bB�����6��(�7����%�[*�+*
�3��y��w��������T�!��R�Y;8 U������@��2����r7�(Y�8{N�C�J��|�\)���|��r��@�;w�O߭*\�o�`���뇵pݏ��f��As�AG��ts�%A�ؽG�ls1#p�T���U\uJ��NA�q�#����F�%$=�s�ԳL�e�yj��}ϼ�	���+~���*2��&�����0�Da8!^��Q��deJ��N����^�́<O��8!^�5��z����l��J��<D3����b���Q}Q�?�V��p�r����TY^j��GMb��L_�H�.y�W
����������ίX}K��Fh���~�iY�G�5�JU7O�\n�U���y����m?ޜw-��t���gռ{j��z��D| 
}�E������?��}тz�R�z81r/��E�iua�#����,����Q��C��al#�t�pf�ʲ��fH�o�T��He�6���u����V ��͘��?��d��䥧Bb��Ŝ,�q��%�{98zc�6IS(��|��y3k�	���a6*d�h�[���?e�"�^ٙк�>���	�oQ�����1�>��UB�V)�at�^��6j�����M�H ��ǯ_�z�[��4�D�#_���)�o߮�NOI@������t��M��X����o:��r���ِ�%]�k���AVK�-����0���� H�� �8���+W�V�f���N{x�0�L�#������0P��	,��N �e?��ྊ�g�Ϟ=�q���8��G!w�����I�E(|���[g���={r��)���,���w���\_k��7�`+,P<�w�i-��'\Sܶ��f�-lj�x�, ����3Zk��
ª(���&��  y�91������ə�:�������YI�Wf9#���(&�Ñ���-�������,������TW��sA���BV���j����Y�lb��Z=��z[x2�-��0⛍OL�^�O
��x�ЖO���~=����/�O�ug��d/C%555�}���r����tQ���������ş�K^Cj�p�{�D �Z\�=��p�ے�/|P���:׿le3��:++uF2�~�*���|�27���g�n@��kjjj�ǨϮ�hV��*���B������h�,��mu��	[j�k��U�D� ��J�]�U��!�F��2���f(���q`����<@���ē��*�cؗ��|�$[Mw��.�m8��~��_�� 1e�7�^�]֘�W�o�H�I\8y�	uqB�.��g����q�"1�Y}ܱ��cZ�m9b�G oɛ~_�b!q�y���?敔�Lb*��$������Xx��e���΁�(��@�����T������Wrc9����\915-ӎ�e�H�o=1�ص�h?�;���5��MO������M����Ғk�}0s5{������,�i�Vyb���Ų)��#��q��5F�	j	 �'��b�\�؏��|��3c}��[=�B	(.:/d0��3c�T�I���,j[�M-�oߔ����ɲ�9WO�BvK[��<�O&t��0;T�"���o�KX��073��� ��HD`���^����іt�ng���۝�[� �gq�	:}���-��Ӹ���mhag�%0_cM�r�0����v	(�ի:R̲�]��y@f�[��~��e�:�o:\���I.{���'�#ϋ����R�z� ~�ណf�tcVl^�-}�>zXv��I����k�����2�[�٣$ ��lL&���Y8�oWwx�P���@�$#�e�Lw��S�ONn�{������
�~�ؘނԋF��Q��qi��J���_*_�a���?�z|���3�#Mf��3��F7a��^ �-����`�^��/���U-��Κ:M�N�S��5�
�	���,���wCFD�NN�ڐ�����M����y�+9���`�-"b���� V���;ל<y��l_=z���-!9�c�0��B�[o�7J���w��D��,��r�:n��yͷ�(�t:u����S�C~9��������*��.�t�Q
�{ܔ��{ZQ4�5`A�H.�,�z���,5]�Qk�+G�s�F�Re�4���tJkoo���ˏ۲�m�)ԘP�ݦMpH� Pp�,=��E����m%��7t~�t�Sٮf�,vD��u� حPBBB����Ø: ���S���.@2�"omD��H���i��s4����~���֩=�ϟ���3I"*2`>�f��g�v6[��
�Fb`�)���1�I`m�v�HT�~�)�d=gP���2/3C���������b9>�C�!gtM�|�!o��]����n}9��*�a&���Do��a��ƌ���`>�0���l]v��[��A�W��`�_^!y��G;�|���ʞ����8���k	�*IU*׳����Flz�)�)�X�"���^<}����h�5�F��܆r%3q��&iǝu�OX�p�g
q� ��1y�I�J=��
����S���&�� <LLL��d#��#��Qmb��`O;�s��(�ww��]Xr�s��� �"yAݩ�H[[�s)F�S�
,C .��.��1��|�?�S�ؽ	PY����P�vQ��g�[0�p���v������'�T����3@7����R����~���55��+�7fy�����=�Ĕ���>�עG7���p��#@7�n1t~	RlT?�BQ*@����a���o�3���#��_�>o��tᵶ��2�"�6�c<^å�5�:���;�;�W����[�T� �z��ʺ��ȧO���-x��,��Ɵx蹫�?�}�,��T���)��s���l�디2�p�2Ӕ0��h_����>��ӊm(�i��{����\�,���'c�m.Z
S��а��>t^�9�ob�R���gq��;�M#9�UO˃s���=�q&l��tY���:���5e�ɣ����d�>�K\L,3,#vx#��X�U�#{�#�j��_�eR~��;�13���d�v�:��;f�{ǟSe`�q ����e���ſ�u� �ϥm������/��T��ԯ�2]@�������_U��fK�l�����*��Č�����kiI���;�@6���4��v�!w�=[�A���@���,/�rǲ�߭�c���Y�$8�@c�T�M��� �>Le)��uVy��f�CS�Z�5� ��Gf�9�,w0�w�=%iQ�1/��Gq��`���b�3g�:q�� ��e�2_��zu��K�n��΀��S��G���q�FMM��9'����ܽ��u:ܘiG]h?��0րO�Z�G`"(�!B�� �8�\�Shˉ^��D��&��̲���J�
+���]�ɧ���F{q�,�����p9KUCc��Ȏ�Ckg[�I���{�>[P-��+`�r�(GbG���..$�\�Ӳ�q�0e��sN� ��|U�l7@���՟ťW �6]��#%�s�|�=��=�iZ�Çuyz#���kHf,�%�@����#x��3���Mr{�"��:�4}}���Ȓ0��vt��>Լۏ�N�+�u�n�w�wc	�~�&�즊��P��� �Q�� �.*�{��J�9�?�_y:�H}�>o��C,�`����>��gqWu%e�z�o	�VYb������Kf��?�Rsv��*�5|�����dz���RG	���#vܠQݵkÝ��@}��
N��UY"(�΢�"+t'�y�Q�����y�u��,���wSW��s����N��n[�E�8�l�<�s��)-�>4J��0��{mO`eo߿�E��(�2H"C�D��z\3Ѹ��c������[����˻'���>q��V#�(t	}�Ķ�������{�aN�$?Z�x
u8����7&�J���f5��o�b`|sY_���-|���)�?�ݻ�r����YA�ۗ���v D���H�UgM��6��oK昦���Y��Ad��E!Y�#t�������KARu�����],�2���Y+�0��E�\�����S�f�2̣�aR�i}��A �nReR��E�K�����L��q���-��ãV�Qk>K�g<�4 >��.�?���E���蕩�W�\���啠,t�����P.I��;v�{�^�z:9���cǏo�CB�+bH��ZF�3%՞��ףĭ۶q����@;���~��b��'(��Ԛ/R���듯O/E�u��u�d$W!v� ��� �����r22���ߘ�ɧ�arC�mt�v	%2vYN��-t��â�G>������J�Y ��ӫ�.:�:Z��nD[����/>Y�>G~,/�}/��d�,����޼yc�/�O?�	�����3U*�Ԅ��y1�?� {ռ���tg��='���(���?�mzQ\�����h�٥v����btt����f����]ǉ������L&�U�
�����Ky���0�23I.�D�C<ـ����kY�Y0�/����3/��Ϗ�v�2��5�Cb�N�ͦ�Ŵ為�U�<O�YJ g��Q�t�Չ+fT�Wc%����z��x`����~~�Kz�f�� ���N�`F�)�ʕC5�l�/�� ���</�YJ�R�N��� 5R��$�"��<�TL����~��.�^�Qe���ڏI�y��+��L}񢢢{��Q����þ�_���U���Ì�ϙ�3ɻ�(���'{E�
�]u1�����α��y3�Bל�K��i^�!j2�*���(�X(S�)���^�_ŧ�,b������4ؔ��O2y~&���o_����S
^-�PK�/;���G�ۙ���;Ӕ.◔��îZ���$��L��6�l������FH�>������}���4ߣ�$���IK��{���gG�-n����^�q蚳T����C����UVT���Z�ٟL��}��;|?��3{֚]D�$Cܗu͓-��ĥ����7}��.N�G���DR;Li}�R�nc�bhfPsС,�G�~y$�=H��_^�6�Q��GJ�wg��S���FX`�sf��z�����#�}}}��G��O-6oA F�֖ �ΐ���8��c��zG9U~U��r�O��A���e`<�*��4�	^��=Ǩu�X�]��@������a��_���h�t.��]�~}֡7z6K<8��T�	[MNٝy�l�:�nSqz���l�:T�MdCW!��`���v�_�̨��d�9�ܙ�ְ@qL_� @�;�SyP�+�9��C=z���n�w.�r�����~� ���{g.��uW8ci	pN�z؃엡yNL�d�E"�/�J���7��#�z6Hf�/a����8QRRR����>�	�}��fE��C�ߟӍ��~�"�I9T����ܩQ�E��`d�
�+'��TX�v��(���R7��@���f8�#�+7 {(��k�^��2e^���!��ݪ**v��^���3���>7���z˪�bM�o������p�Rh��I��D�Z��Q+n7	�^��Wv|+�Ԓ,`o�[lGg�H6�Zܮ�U��1�O��2�-5�A�^F�ϞC���V��?�vpx�H<��͢!tŘ�ڣ�F����W�p��3 W��5�Y^_N�~�s���jQ���}~l�U���Q�ɓ'��atSŠY�j�9;n�*i�l�O��:�EpWe�����,ҟ��iِGΗ�L���Y��w���j�`��d�֦R�E���
���cF�2ؼ�СC�߇�����U{���,ӝS�c�y9b��M
mj,˦�����7+6��F����x7
�u�x$���o���T���|�m���I��q��C�N����(u��6;�X��QV�E����8B�n��-!w�u�)+�:������g>��¿h�>��EǇ�j�˒��U`
�i���.*����mUG�m��i�l�k����ڮ����}( ^�;O��d}�����񱂪trc��.�ըՆG@6T�.(Ne;34N�M����%ٞ��D��P.}
���[1;�/:z����Y���	�!
.Z_��$����A���xl�n:ai��,@��>�9���0£=)�6�*����b�d�}�9���eg/� ߼e�`���X�X���(���a,��r�؁����&�y��Yڐ�b�~�<��l��w{���3�ǔ���<̀��:��;���H�9�y�D�Mw��&
];]�7 +Il�/\��q��+�`�BAA�e�6�]�2~w�����Z����W!�73�2��nd����������"+#��p�����D��� �?�Td�=�_���jf�Mt��������u�(�1�,��P��&4�H/]�j��fD��}+'���#����k���ﾠ��N����������7��|f�̀}C���z�����ܼ�Q�D:k�f �qG��hN�ympV�0�$��)#(��J����`���U�����####���Z�1�t�/�l�UN��}VUA�<H�+%P�9a��_@0~�	���� �08�n8�d�3bU�I��o6;��i�#c��!���6�e�p.��ݩn飠�Qھ? H��9���d��.,��0f��`���N�BAY��;_�4�|]�]��E����HG:�Wt���}T�>>8Ш���+�R}&��G,�z�^�w�,�;���Л�����6��3
�w�
���qAzP��q�6���w1P]�b��-w���s,|v����x��+��ЁR0�%q�߆��=���}�1F�/� �����wO�m(-�����%�2!�<�u�u���7��P��[���F\?�'?���C�}�F6Nk��jȳ����'8q�{?ٲ��l�ߌ'�k�|d��nO�����;B�)����ӥ�k	*��Ag���y�܌b��XR�Q��1��/��zPR���HG^�sJ��� �{N}W�-�c��CڤK�`�:���'"�4m:����8�^x�����5�[�/HN��b�Pa�)T��l{�(NRSl���0������+#)��߽�m��m�j��U%yJ���{��>�2!4��ɣ���&}��b���%��m1s��Y�})Xɡ<�l��(��ҏ��z���s��|xs�z5������f�"���;��Z�������\,�=>3[��Ӏ�%W�Z�����4F�����l�0���,��E�(nZ���R[�����d|5���_'��s�A���e�ctOa�����~�D�����B[@L8���){��k=`cQ�XӼ$%�z�C�N�4*�Ǐ-8�S�TP���o~*�J1�zZ��Ѕ���l{�ʭPqypk�q-���և���o|d�U2pF�������EHr���kQJ?#SL:܍@8����?��? �y�9l������Q��K7�2w2��JWzv3��׃zr�OZúm�����N�jԃ��r��j���B �k�3JhT�i&���`��5�;���]�1D������8{Ʌ�&̈́�7@h����K���L��1dK��>Hހ�fC���H낒6���?�h��f�R=�Y�?j���}~V-"��ڶ�^6�Kt?�Y�ϼz���Qz)e���NmP��j��#��C����bR�9��j �4A�m�=L= u���X�S����̚�XS6L�(-y^%�`�C�����\��c�9�4��2M�0�2{%^�O���7��=P�?�����g��wp���;����<��IZ᫱%�5��-a>y��G���/�"Ua~�G*.�y���}$������ZUŒb%��/��3	\p���۪2���BZ�O�Ti-�K�zp=g�a��D;b�#/r����'�K?�p�3��������v~�W�
�z�螚(ʤ �(.ku����aĆ6�Y�hմ�I_��B�y�<���:,*~Lo��-J�qJ����_<����~�翥ݺM�F���5�8J�Œ��3a-������zE�HpV����)V"�p�e�Ѻ3<��Vn�Nwq�2����[�����WH �n�*��eՑ.I�͝=����#n^:����M>�6��U�t%�ƍq�$��g��L8<xB/�{=M��)�}g�Z��_2N>ԥek2��-䙊A(2h��]���sd$#7�}�������6"�Px4h��T"�S} ���=�V"�S��rO��������������8�ƍ�?)H����o>AxR$������l���7�ꓘs���B�&�[vy�'v��Å�Q]բ�Z�5`�:�W�GJ�2�f���1��[
,��������m������n��'��o�%US����#�(Z<ead���JڭB����YrcE���eKH�^s�\�8�5�����N�le�j������o����X��J�'�.E��(,-'���裨�K���*���S��裞YO���4�E��q ���e�L�Y,�s�)�������,�����Kg�Zr�*3��T���k����2%�(�悫m��]n𱹺
N�;�%7��."U ��+��A�1���%?))�J���ND|�#��������YdT��b�X�Lv�"�)fϧ3u}}~������	���g�hk�it�{�	�,ħ~���m����sX�w'�}���m�bS�O�߉>+�q��#:�ن:��V�y����uZ�v���)ی�)���U~�ZL����vxBp���L�n���2�*'k�ӈ��$u_$����_��kgØ�5�g��o}h�Q����z5<F�%��ٿ�::���EFF�p�����3�K�č�;Q��Ҏ���}�66sB�$����/�xa�ev����Y��~�A� Y]m�V0�L���a��|uP(�o�����=�\��Vo�Y��)ai��z����>�-���R��~��V�zX���b��P�?���s��]WP�� �S-X&�7�C�c�ћ=�8�W�ldݷ��K^�QĪ�s��w���K�l�e����tY�R6<�߆�Y?����vvv��@���Fܯ�ϋ�Gm2���Y;,S�t��-e�`|������4���������W�u&��A���߼_���߰�8k��s4��(�p��k�6�^���H�Ք��v�]����/C&Y�B�KG��~ry�M 0V,�P�:"bS@�	�k*33�2�5/�I.گt��o2�rz��x�ʽ+/hy��*�����P��"6��
K!zw��*ɼiǉ��b٣��K�zۊvN�ɱb�	\cӳ���i%$i��ɄW��L�U^�`OS��`C�/
EԊ2��X�z�o�>��%+'�<����)b>eCL��6!9�uC��Nn���#|��e��H�I�9O�}>MM����ʢ�����e�|#b�u��J�r���u_DC�+�XQʩ����
+N屢^%(���`1�����n7��|�浄]���~�AY�7�K#G�u������N������t�GO"/��䃣ӦFK
6p�}�0��Is(�ײ�����[^<���I���y�����}ݛȓU�AS���H�he$����/B�[1�lg���a�-`�m��5��d:L8a�Uq�vk@񹡣��I����^!��=�d��'"ֱo�I~�?�J�NY��:Sz�A��%����|j8������E��;��v�3$���kvʎޏ
�$��)Z?a�๙QBU�nZ�"��$%,Ri->Y�U}:��4c:�X�D��9?�s�VA��,v.�$�O��a�C�#;5�_ 8, ��W���׭lDs���A5���H��^P�_��3b�(Z�����
^ş�so�FQδ��|Y$��YxOe���\O��:��䢬z ޙ����W�w
�u�q�&9lD���m�\pE�����!�8���@���Լǩ��d����QsCRQI���g��q�/���o� ����l��
 ����^ �n��Mi��~�bL�'�;y?č���~i����E��IL��{���Dކ|�5p�Dd}��¼��ln�'���BuYŨ��i���l����_��(�� �Zp��3�`y�K�(�S��n>�\�kG���oh�oؠ`��e�b�վ�ph�`��߰��L���o����X�!3c�ӻmQN� jg�w@�O����6)�O�ۤ5�������s��z�o�\F�p
2*�G�xbA񎼼��K�}$lc�"=�,�D������ؓ�4�1y
{��4@H�:��j��We8v����sx��Bt�\W�C7� �s(�S�`=+Xs=ĩ�*�RΤ�A�>� �(#��u�wqr`�\���(y7q�2>�{z�������p���B'ʹ&����km��o.��fT�###.�|���������D��pG��<.��s,]��c������ڭ����L�xw�R?�DI���7E�a�= ��8�<�F�q�"ll�7�.�PL`3M�9'}T�4���	W^���21J��U{�6zƍ2���Jէ�y������D��{�<��z�a¸
�P�*q �j.l�;����W�m���J͑�:s��i�u�"�=�
�@{E�:5���w�|kln ��˾�5�<����)�h��<��R��x��i�����'�B�#>���З.X]�
o���l޺J�z�榠�1g>����;��i� Bu]n&�C� �T"m(/�°��T��J��a��0uX�
 �w+�B�Ve�=SуH��j���{�v��]��$��&G����S�<��s{��Y3��`뀦"��=�W�ɻ	���N�"��b0w�V�ֵUR�����Gv,�	�m�8*�%~���4u\ƃcw�o���5u�<��+�N�=H"�bI���ꭴ'VP�����^`eO�g�E��]�@��p����������H�#��v%!@2�8}X�����Z ����[*d;���o�ğ�ރ���3�]{��s�c�������V����3��1�䍒�Wo}�`�m��	A9>���ޟ3�����iU������%Ho/	�)"��8�N}ga��W���:��خC5Fԍ�^�Z��1OѰ+���ltv�W3y:w��j8�!A(���K(�u�U���k��/5c����7�KЏ	�]��V�F�
�sv~7qj�
I�XSSL��rl=RqԤ(�p�����lt�
]�����_l����遮�����a68�E~s�-���h��6S��i� ^Ѣ9"�(/�D��D�����K�����z��Bc&��|�5��t6�!�Z���$o�
O]USW���ӛl6��ݛ@t���$��!��(�ak��:͒�ӧ-�~��i�|'96��w�����{�e�u�.���)i}[բG�]�e�����Gu�N��d����`2��=;3Y�"��WÍ��kT���ύ��w����[x���"2_�b�ҏ�AE�yk͘����{�5�,F҄��㠖*;2:*)�oW�3��Gi�=�!TtZ��Q*���R���Yŕ�a�˸�Q$���eZA�w��U�!���@E|�LT���zB(ۜ=��%ɷ7?�ue5XΌ�~�9�������\�ʺs�F{0�z>�T������b|�����1*�O�HԶi��|�i��p��,P�ux
׼�K(/���wSْ�G�#�����7�9��hg���Ls�0v��a�+�r�����H^b�� ���!n<��1Y � �⸀/Vn��oB��K�Jg#�,��$� �C+p3��U��bX9�2�b��Zۋ�`
V	-rt$yQ6H[���C���5&�d�z���`:� D���8����[�:��[���!�������z(�9<s�B[�K�(�Q�X�.��33�$c�mb��aU6������F�*�p�Zl�!�Z�i�E²"c�J:^��"E'�݌������(�'�)�Ʀ�8��(֌E ƭ��U���1|�C��M4U֭;b�'��pQ���/�5v��2Ut�w6o �_%57�8.0��SI ??W��,'�Tm���Q�E�����:�l4���_	{�����H#�U�5��"%�x��`�ɯ��F&�{0 ���P���$9�s���K�*|����د<���H |�c�[�Cl)o)g�8��b��>�v�-(͓�U;+�-^�j�6�MS�g�V���A��^��Y�6C�v�B ����l������׵��=,k*--�RC�t��Ll���QIR:��4f�:P�I�D!:׌��JB�j�Z�)�����yg�����o��w�Ͼ��^׷5�<s?������C�s���sb "t���_a'b݊>#���ޗ �ry��hmf�ZLc������ԥ	�e����綶�gQ��rY�R
� ��+��ÞE���A�@���x�L��vݳ˿���>������i���ɕ����_K?��?S��|�&kN�4�Τ��b��k����_Z�K�>8������Ώ��`w�jd�hi�? r�ic�i���Q�+��H�>� ђۭzQ3T��^	����rb8lh�T��zC��-��Q��_���'|2����ь)�A"�7�O��Du���７�gt~��Wю�G�=�+�*0f��V�K��*ҍdo@��m�����|D���K�ws�d�%]�ZG��&�c	�"gk޲(�4�[h7ۈ0%��C��ĿJ�?�G����?��𣞏���� ������i!K�^�x'�Ek��iԎ�s$8��~ĿnF��k�������;��6E<	,��W/�e?�+����a�~���'���eq�^G�1�̤왣��g��8�,��}1]��?�h�q��\"����/DM����z6h�)��%� R�i� �ۓ��8���W�����u�^���]z�N�6b;�b���y���;��ź�Q��S<��s�co~�21\�?�6C�S�u8v	g�ۍgQ�;�O��:��ٮ��J���3=SK��o�4^<�݁�����cAxqg�\���-�����!c����_�M<pq��H>aQr�q�ϑ�hy���̳�9�_!z�$�/yz2�_p�Ox�m����_�M6��|�3�_z�=wk܋���pC���QY�
���ˢ��]�l:&��Yׅ��~�P����N���`cy��W���>Ӏr��4�����W���F8LS�+�,��b损�y-�D,s�kb"Q�$׶�rY�d��X���gj�R1���܏w��~��}�LQb��ecy��i�g����|�g-��v�3���-�EDK�ю0�]���X���|f),�\ԑ���vΑ���� qBe�Tv�~�M߰�M��0����]z�k��,(�a�������v�x8�/)å��[�Qe-p���uy�����3�Q�?3#���
�_���f1���a�!�#���ov�����_�֍b�ܗ0)�1F��.��X���3��]I?& ����73�#AFr@�XӃ�~�G=�ÖO��dǚ�B`�'�� ���\��;�mj_zV��،��h`w�Ư��7~�0ش Y�%���V��b!�8䇲�=�l�ǌ,ZV�跶�&���}�=5�m���QrϜ#���fQV�#�ٲ�3�� 4F���&��]���}��3�0�w7��̵�.���|�����T�S���?�;t�;Je?��w:,�W�Ա�q��Z	�|��7+���8~�'3�vVb�:\�61�����56��}gV�����ݨs����
�'�qٔv>��G{f-�bU,L���&e1+e�y����,��:�b/�W��5/��Ȅ���6J�c����n���|�c}C�щحv�7�n�1~�v�S|�<~w�������-�v�� PY7*�0����$4�ڮ��O�uj�㯲/(��>��s���	����Ʋg}�~ި�fC�}�9���P���X��.���+� �A������׫	J�k�Ϊ��б�
�1+�g&��"u�O%�Q���j��Ǿ��
����c��� !���b�F)pI�-��ج����s�|�v�[�6L=��>��	���k[�Yuy3���U����)�۔R��O�:S���&��?�.��˽#]�(���80P���;F9�"V�{3��B���cqՊ���5�w���e���^�t�8wzA&:�ª͙�/���C�+�0��m�Q��^����b��]E���F�u���HI�P�)�����WJ/!7�-Xv'��$$Dٝmz��u��R����!}{O��F鱗{��̗�)��2���'ގ�����Ѩ��ca�#X]����5j+��GrEN~�l�ɿ��N��0ر-L�������H�����xt^wR��0 �I[�vgl���_%��l;���`~Z�x�C��=�N>�����<�!���x�'����~�������	�stb^R��H/�g �G����U���	xV��{���DY5G�L�D+w�I�lK��[LC�h�c-"F������_\�y=|�����2$_�Ѩ�;=�%h�a�k�1����E+X!�����ǯ
S���T^��}�鉨��-s&��۪�LL$`k�����'0�j�'�����0<�*~�W�Z�����Ic"��%�"�(ռa�,�w[w��h�ڮ�ȍIX;���A�[x�����٪)fѯ���3��q`4��b��R<ğep��{��*���78��mw�nhx��X�[�x���f���'����ۡ2���b_��2ib�Q*8e�O��\
���ia�;\BH^p	Ib��wl}�
w�e�"��&-5�	��`<\Ҹ/��Vq�i���:�������Ɲ^�A-��|=无��^e�R
� �];����q�.�P̕�iz���Wz���:6�`�9}c�u1�(��a�RJ�L������)�!�/�����[�Gb��i ��n��q)5����,�2,g�&����9'y�~���W�<���{CK��U�CJl���	�\pq�ֈ��jo{g�q�L��˸2�~�.��K/��j�|r4UQ.V;-�������ӎ"�_^+���t�ݚ�c2�&ȍ��xˉ�n} ��^�_&���NhZ��k�/�X�GUk+h"dM�}c��e��<��"�\D1%5��`�"<�%W5��-����	�;O?�ͨ枞��= �-пϫ��aҒ�Ol�i$��U�-��1�D�x�f�'��_��MaD)�
r���7�0AB����Լ�]e4<쐴�4���G�����9_r�Ӡ(tT��ŵm����� z����z{�8�щzeL��� ���i�]�������A�m��1���J��̚p�k�����٦��_�=�O�+�����Ǉ��,�G��JGS9&������X|���~fk����]�7����e�P��oE�����3��Ϳ�G��LP��̖�l�][��O7i�Ai����I�ԅBs��`��%��}f�RyJ1r��vi,X~]�fL>���Z�¸��,���اYP��E�J��0	q4j)ո�#���(D3"3������s���-jt�Z�x�غ�X$��q϶X-�R��Yr���:ʬ���>��10xR�O�H�^��1h?Y,�x4B����U�yvzI�┚��1^��<PY8z! �&-yU�0C*���I|�w;K͡%�9ֹDk��B5���D�V̼�����	QCM�:��)��i�n�2S�ro��#�s�������Xi��	�k�����q����)cDw�7H�/k�{��ٓ���qM����� j��V�iip@��*��сMh*s?_TE�MFm۹�]�[Nn��Cs�a�y/N�p��<�l����|Y.�ɎۢD�3i�CB�(���T%.<W��Tx�\ݵ�ZX"����o����[9:�z���.myp[��:�����T�G& ��v)�n�W��}pG� ����F�`Yx:q�f���7_���F�]74$}N�^7�XǒOx�A���s�c�*�/��r>;&3�i�df�����]��hţ'n�r���)ɗ�W�Ae�`���?X�{˧��h^k�Z|yy6O��9�iW?��xI-q� #�kAw�XT_��_���q�ĺ�ʱ��/�bp��Ґ�<��F���i��:=7�{�R������EW�io��/şsCל�����<b��8u0C9�s�Hz��??14\�K�	��)s��)b��B��6�3�.|ܱ0(9C���8��E�x�w�>��]A �_�Y2;�f��^d5#z�$a�����qw�����l]��a�5�\��S+����-]�
�І��5��*%�5K�h�l`��;��-֢���Fb�fԹvM�C"y 4��G��#�9c@J�G��j��SL�)D㑰��"NJ��qH�I"�:�˒������P"�����k��,���A岡���4��~;�s��"�e":� b�x������{o��1�ba3�_cҢ��g Z��K�5���P��[�v�z|Ӊ��M1����8O��0S��="K�lb��q�y1�,������/�2����R��x����A��B���C��5�+�Ǥ�^	*/� �|%�W��U�\�nz?���)6^�����j�D�K�.3�������J)Q�O����v���i��#6�ר�h�q!���<�Ǯ�k+h:��מ_y6�93�vօ����^s�3Zy^�aܬ�?)\��K�OG]4�M�Oms����Ǌ��ĵ}C��T�x��Ͽ&-����|��{�kw���n`�*hnYe��RTGգ�<O�3�_n��-I��I���^9�J�{��A�$��v��G�s�.����79���)T\m�l}��v��aV�C��Ŏ����s�R�}
;�[��k1��
����}�J���\��Zۡ�{����O?�Z�J	6kYo8�v�\�D��>gRc�+(�#)&��G�C��Dl�[����lH'�z#�ӺQ�浽�>���A��{�c�癘"��5�©��w�1�!
���X$r��H:i���^�){����r�l�󀇱���_�x�v�Jz�u�E�H/�ċ{rMY��&61�ԅ�����+j���@�"b�\��keu�)~z�3�^�ry�K�Ӿ��O�Ȇ��Qh�i�I�����l�Ǟ6eV������L������<#��*�bZZ)5�;q���s1�NN�9��{@�ss
a�R('��޴s�
�:���n�l�AI�>�[Nc|?�ZSX:�����7Jv�Dr����������,y��^����)=^�ܥ��BW���Cc��a��m�~۝���NM���0�2	�%Q��ÜbU[�u�4�;��5�֖���._n]�%kT;m�h��cu �S�mA�Pi��$.�2]�\�U�Ph��!PJǉ�*67DlU#+Sb��`����aj�e��<�@e�5�|�q�J\�$c�&;l���-��J�|� �\j]�^��~'�"�y`G���s�����L_~ݜ�ꦼϙ�z�+N�͌�i��?�B�m5N��n��d�s	O�\�[ns��^�M,�R�M�l������^�}��ўc,-߽�|%��'B͏������z3ţw�"�^���w})b���u�.�ig҂سհ���'bsY�НF��YJ(T�!.1��;L�k�8V*l������~��������q'���z�� ww�b�zaW��x$g����ӎ���n�|�10q�5��=� "�7�c�F��P��?���7�G]�x��1�wlQ�R���U��Le�T�r�����mԜ)�DU�O��j��D��"]�������L�i�$�5;�m
Ϗ�A���a' {�x!&6����	��I�(O����a�Ӛ9o�a����%"Bg�ڻ���oʻW�*��~�_�4�8Ɉ�Oܿ=X]a�db�m��,I�V��"�*���'��X��k���|�z�M��J����$/:}t��ܽ�q4�Jcz�δP�١���?��	X��	/f.�n����n����Cwc˹֍�<�x�#~��"��i��V��iҒ
�����c����d��?u�� ����^���A�a�>`ӷ�����,Iፍ�=m�ð�TO��3�'�eB�_|�����Q���Twz�a'ql�G��f�����I�܀�'�Rxڙ��t�y�I��}f�^�3��ojV� �1'�y'�� �-��%�����ϖ��z�v��)���)�?��Fb�֫V"�˒�lJ!���������~C޶��`�!������X(&������Rw0�=��9x���#�"��$2n�6��`�<_ B��@�\�~��B��϶�t������"9ǞR�@r�2'����Փ�����NIy�܀�݈Cx�;��,��>�Z1��h�824�����5�|�Sb[���ii�zi������7���>ifp/B��ޱb���|K�g=�ܰV񲴼���������6�{T��Æ�"���3��͗�_@�E�Mjz�]�z*�QS�x�8�Mw��/��N��E���OY��]R��Gr����	[�|��
&��}�����$|��o��ym��MZ2���������^�Zx���V+��ޚ��-a(i����%��Yc�m��/�,֛8͐��w�hl��^/E�B#+/�f쳼�=O�ms��ѳ\[:�Ķ�-��EV�e�=��M9���q�g�h���Ϡ�'�nw�U�cʘ_��݊����x\Z�S	�.�����w��}�k��t���]k�g����)�A�b�7�Ǆ��ZOd�|�$lVJ�Px3��Z��*nY������+\�Fb�`H�����c��ܩu���&ƢA5X\�
���	�ԍ����8r��A0�m;�:NMq�����$&(���4����ĺ��A0��>I5��
�ޓ�͟�����w�R�j�2��-}v�loIX���Aq��L� Q�t�@a���2�O��|K9fɆ�\?`a��1o��'�_,�_�����VOs���2a䘙j;S�m��J�n]�zh�+�q�n�痩�J�D�D+� ��lQr�u�}�H��3����T}�k��ﻔRXǃ���V$b�+]FRS����yu�/:bd�=p��`|z��,�:3P�x�u����
oSF3Z?��n�%�G׏�_*�Ë��Y�������؎����<j�E�&x���i����D��a ���-#�W{���#S�����L4��LZZ��k�$6"�j۰T�E+���}z���s��a{^��&g�IK+dN]ڈD�#��RK��p۳�ӑ:.���Tu�%]j��־(��8��[����͑��QRU��j�p��f�ٱ;*��	�g��	�,6�o;p?���π�� �����;x;����������O2�V����;��ZiҢSjj��[�5v��ы>��-km U\|	!{�tզ�J��)��O% ���5�o7�HD�l���7>퀁��%2����-�y��A��<ަ'�/>W���y��f�$�3��'����z�_^�t_�W{�����ۃ����`���w�8�(ݭ��x?�xu�ppݼc��R��x�7w���u^���@�����Du�NİVc?�6n�(xF�-���c�u�V��k���!E����dxy{P��ߵ��H/@���y
�����4��I	�����1P��`��"<����y�j���i���Ay-!�wp�S�݄�Xd�Ee�뵱ç"9�O)
0�4�USJSxˤ�����vu�BF+L0�t�0�WT�%���L�{ё��!;R�iZ��VE�6��i����h���SS�Z�֛F�m���$ę��η
e���qX��J�T����	99Q��&�|���R������f��͎�����C��L��7�?�[J�*6�R�"A|�0װ�4�*�s��6��EJOEi�� q����F���M.�����gJ�{�ji�1��I6XZu���Ti܎�֮NR��$���f䏆"�����1J<�np�&gR�����Pkp�E�Ə��x\�'5.ˋ����H�)Kp\z7�Di0	�J �qí����XʰHd���Ϫ]{A6��=N{.�:�y�ӽ�[��*�3q�d��~Yt�t[��4��<�t����Ԧ��W �Y���T�ǻ3ܒ��MTEMIjuKg�B����,�dɭ�k6��/ٙU!j��H�)ɋ�A�C��K;���v��[�*�GJP��4$¯VJA��,xy���~7K=ֹ �UV� ʚ�)��:�����$�s�&��i���|��>z�|����Jw�v��`�!�Oaխݵ,!7�&D���]C ǨΰR�?)�ф� �J0=N��F��##��C����B0�{�b/ɤ% �` /�B��y��|$����6���Og���b����X�F�ܫ4���Ir:���%�G�.U{$9�B�#��S)�Y3M�dV��*��WJq?4^��{ْ.�e������(���^�+���6�Ȉ���!1�d�p��Q�<W=�s͠��Ep(����Uy4�2�6�w����2����}rQx^t�����R{���@_�○�Ƶ����y�":a�<��������l2
�v�oPoݶ��ߙǾ�2��T7�jp�R�5Y���Fr�`
����&$$��qa��U�_ �#���ʯ�b>�?����.Ze��}�:U�7��A�9�S1��=����:1�C�-(���m�[	�@���]�1��#���<�am�^lZ�5��w&�	�Ǌ5N�0 et��cu�o\�2� �е*wg �i�ZW[�J��Ϥ�t�E<�k�	P80�p�z�,�v�G"��"Z�Ҵ��q]��@U՚Lw�i�/'ii�TU40�Z��!1u�wi�wYZ�DH<��,(��� ���d%�h?e���U�,%lp����QcR`�^ �]�F� Vw����$Y��V�L�Y LЎ�a.ht@�2c����?�����+�㺺/Q�X9j~�Q��Z�H��ۍ�V��5�Zj�nX�D1��x�<�(��ӘǗ5�mp�zef�bj�R
�.��z͓���jhs� گ��˒l�Zg<���FE ��$��1L�5R(|�3(�ſt�ʹ���q�!7�ħ��s�W��wm;�b����,1�)�U�XZd$����K��W_���7S<B�SE�7g��U\�}�y���I�ފ��C�њ�6wbO���@;�1?E���֕�;�3q0?h�/C���)e6�����^�e҇5��pΉ��j&�3S�6BRE��\��Tڪ�L�ʅ��(ش�G���J�G(���ށ�(DxF��k+�c���1����(�*U፬d�>x�fR�DDh�b�j�@��`sr�\�~��Bo����ٲ=�OL��j�n��,H��y�V�ӱa64���r+�*��#j[���-�6{�KtdÂ�A�s���y��
J�m��q��m��!����}?�Գm�dgN�S������J��Q;���j<��+a[ �z[�>	��t���A�-�Sa:ٚ�;<�i��M���4~� '{��If[q�j��ش�%�)!.u���5���]R+7 ���j�Y�tA�vbM���(&�.��~��"+�)SB�ÿt��q:�C];>-���c���y�WW��Ni0�N ��žq8r�Eh���w�vwFLޱ�2�1��VI�.��$*�r\���#_��;�>UO��(�{�0`2>u�m�������z�\��M}���/���7����N�I�h�N<�������6�AV�EW{k(Ȥe[
a�dX���o4����VR� ^c���I�[�+="����Ձ(9$r}�lI�0"9�K���7l�Ǘ�Oj�/$�CP�V��Qfc�%	��ّ�ڇHz�bF�b��S����L�3�$���H����v��xQ��{�����m-��/������$&sy}@
r�]�ezWJQ�J�nN��삧�D�=��gmK6��C8p)hWf�}3i������ I���^ �`��"�sJg2��e�/�I8�u� ���ا�}�����F������f)�ܕo���{b�j�)��lh�QK?��S���B5Ț��n�ܥ�[���� ؀<�}�����7�փ���=���U:���Z���GFr�d���a����
:��E�G,�u�H�����K�z�E��� u��Z�ԳN��*�!WK;��.ź�L@_� �+1f�9A$}~Q���e���)���s�C�7
j�g.qV��B��vEt�������$����=I[s
A�N�iO.q'�W�oȾH~�e`�� ��٘]�*e��{�x�o���k�A�ëݫ`O"�7>ʣL��ھ0px�BuKw'�s�4��S����OI�MOA�VP��[ہ��\��a0m�S��n�'i��e��I���6�h��b��\ǿ���
���Z�]��=�E�e7���赉���S���#}APա��-�g2O�P>H��	�ڬ�!~��N%�QM��(�o��"�s=�SR;�?�[n �8��L�>�$�u���q���T������;:D<2D%�lT�|�9���Wޥ�a���xm�C�h@}���Vtˑzr����V�3r�uw���_t��^�S�B�8��"�;ߋ���P�}VC����un�pV�ݨ�a�Ҥe��-�a��{�ܛUƨ9ysc+:�� c�o;��;�?�
�z�֔aՑ57�A^s��԰�kO���n�/48Q�"vb2{l[�ĮuO)��Ů�{���D�F���pw�Xv�r._n}M���M���KR��]�D�8!ٝHCt�&�e����_�0��z��Ց,_H�Q���잵���GR8�A��4bHx���#@�j���g��jx��;B6%����t�T���j�v��I6
�̎}����w�F>�Fy���=$��9�W�P'z�ɓ^���w`���[������U�z��"�{TJ�E�$�)e�D[�@
�r:@-gǵM����|�$� �:Wa�:\�:��J������<T����~f�Xo8��9�u��kn)�n˼9Q��ĒǛO�>ܴ0u���eNb'h��%�d��f�ɶ�_}��;��vo<$��Z�ԭ-�~�(�&����	�륛򟷬��j���dcfpW<c ÝQ8�Լ�i2V�5�$be:�y4�n��Ǖ9p�-jz9�Ҟ���:y��}4�CUU�?..nxz����'_Lp�bS��e",�t�b4,�ch�8����qv�[2�C�Ө?���N��뵩�+Bq\��FOzf��hCu�-X0�A��jW������i�r;�i3;Umv�(4���_<��8ui��U������U��ԻC��X�~4�=0f?�rgՕ��G�2�z��^Ґ6B��c��4�!׹�E��<�;��ѭ�C�K�&����f�T�rY��ǏmΫ��Du*���������A���{܃��c%��T����=N�Sl�������f����m��\鲝!���:򔜴4�BCw���j�I�����6��rp�W�X�2[��23��o��]����'�MU)�V�:�B���Ɓ�.u�9Gx��,�os0��0t�9�9���aB�<�
D�Jx��J������������	q�w�L���TH=
���}�e�>.�?�RX�kCOϒʦ�u��[un�Un1^�4v�b��$E�v��;���Hvg�E���ڈՖ���w5���^�}�u/�տ�;%�6H���(�]�y�P�V4y!��i߾jW�j a�@��;�P$�υsDD�Ŷ�yW�<RvG�"(�VsL��7�#���������ٿ�R�lk������w����E���:���	�}��E+:C��~�Ԧ�А+�u�9�l�㑋��S/��_��S%�}�HLQ���#P��O>L���U9������p̥�ss�Ɠ,��&-Z�o�كK�,�������R	�A�1�n �Q�;�����L�_��T�wqMp����8{u�
�VR��2����/�)o}�gJ����`�IJ)t�H3{3EJ^	�}��X�������C�W�2�P��~���Ab�����Иx3�V\E�����%�'Zs�yw����fk����})s��B�Oa6r��h7�e�{~=m�q`�K�c|?n]鷅4�{��CC��(9��o)w1=:�uقԞ��5���Jի��SF���^REk�2 ����d��:�����I֫����ty5=[.R&��]��9� Q�&==!t#^�q/S��=y��K�sh��a�1b6N:�P؁�/�!�Zn,��E�9���^�d�Ѽw�m�p$��.������
�E�~bb� ���J��l��	��RLj��H�_����UƊG�R)� `Zl:M@�7�;\M6�HZ�@�d'Y�)��G:x��xC��(��Hz������v�Ç�:�C�D'3STr���T�$Wz��
�_#Vo�a��8>:5>Z��D��M����4h�b��C�9�����"���o}�d�C
�y��ړA0*i�!�
I]�xN��g z�Q{��mu�ۙK��F��,(I�5��c�`��iF͓�i�6��
$1ҽm��Bl_#�C6ZC���(���@��!D�7�p�g�+g���z�,S���k�/�<���Y��[a�T�_���|�ѵ��� oV^b���>�+�t-��qt��VI�4n��ǟ�!DCW~@�Bӝ��Ng��4�Do�8S�9�������~!����mrW�K�����~��ߏ�6�Z�ƚ����e��.Q�����xr���c�;I6��L���U���H�<��э�#;�O�bZ
|�!���}��Lrǜ��P4�Z�ٱdu�����̏��2�֑����if$�i^�
)a�)�Ð�&����=*mT�	Ϡ�=�^�1�%O2]w��Gv�zk��i����@��h�iD-�#خ��J���ۊӢ�["�TE�c-X;�r|+�-�;��u4�[�Ң�h�+��#N����RJ��<(��;�ӡN%�.܀=�@�v�WV�R���M	>�t��
�
q���(O���]�k���_H3|j쥈}M��_J�9k1��o��	P��r:my��q�+�3�	0y���4^�qˉ^���C�n�}�r�9�[QE�z���l�<�h6z�M~$����)��K�M���R c�Q�'�����kj67=��M�.K�`�`A�4�Å�{h��^����&M��8O���׮�[=_��r&l�{�gI{���!����Lq?b"Z ��$�qh�&��M�>Pk)C�^N[@�7���c�����i�x�-��z������vc���)R��<��[ed�� �"�ģ����:��,#f\+\Xw����R�����n�k���h���d�T�y�3h�<{�V?:"���D�}7��g���Z��ƈ�>^����G��u����T�����¸1r*��I��7��H�&Bg6H�)Ǖ�f��{Ux4���-�>�LXZ�KT�ۋ��K���ߒ�9�tP��!D_���E��}��[{��?�w��O�>�Ϙuҧv6,;S�d]�պk����oD$C�`,O�]!�4�����AG�xw��ͤ��%V+��@^�ı�?T�C��c�i`F�P�Zn���Kz��y�kkO����.0'�pEv�R��U��B���3����U#���~�?< ��'�s:�<��pj���e������������bG� 1��y4�'L��_��Ӟ��/�A/	ʉ��"�R�+��;Oix��[H�tV�
�Z�>(�����sZ��:�P3���AS���A�mց�o~_>�"ӣH���g`)�(�&��!
;$��>otnE�6���a��?�̋K��0/N��P�	��G�u���F������A��ǰJ� {�l��Z��q1�ҥ������j3m�.�'�e/C��z�=�-�t���je,��%�J�0����i]o�����oq��x-�઺z�ⓚ,/�v����.�ø*D����χV.� &zm����I��(��4�ԑ�})����4,BB�8�l
G����?yRP�#rU]�Wu����6�+���p��zIW����jMk�I��ǂ��� ��16���B@x�d9x����h(�q��HčN��O�~�t�zA���[���ufy�;������ʦ�7����=��K^=� ��T빉�2���j����Is�h�dB���J�xw|���G9�Z�qmn`9mA���ME9~L�o���V�cU��u�<Zy:���E���V{���ɋ0ۨ��i�p�?��<c��rA������7��J�������:h+�G�[��ɪ����?~�n�ΦL���/�������+�"i r����H�p��Te��!(��xz����d���w�m���]�u4�v��ȕ�W�0�`fk�/�h�^U�kh�>�Ⱦ����/\�ؗ��;��8��|�E'On����<���Gց�q�z!�2�0�����Ե�Wſ�#��l#��BV�
����S�Nuo��y�K�.����՜��}�n�vo�}�C=�8С:,-�	냶5���Y�- ��%x�3�r��A�#�zW/�S�2������wZ�؛��Ke4�v���P���_�I��a�3P��M��]��i 灒��s�
�-YD���A�7�S.�����y��&��S�j��'�
q{���7#�*��;=a4S����Y,�s_eNpD���-��f#zH(�o�b~��z3�±�nŸ�b���������Ǧ�����)�[>�ۋ?��{��rb�2f6ɪw�x�	��=\T�\&����(&�p V����Q\o_�4������e�^�����B�����Qn���V�Lz�(���6)���(��+��zb5+�Z[*u�h�߷�R£�_��^�vF������I!��
!�C��.����/?��y��ˏ��mZ��� ���'��s��*uɍ:7فφ|��![���4����"�LS=���5G�I���L��"�]��L`��;�:��K	�������[���'��|
Am�u��caJl�@g��f�)��)�[v~R������^GAn6���&byA��ݘ��sk��}|�1���b��	w�UM�)s�kQ�y�BH�h~d˝Y��5:WA����'���jPN����1�@���� ����;oY1��@iAzP�-z?f���OK+�V�{�n	hrP;R�M:���&��w�ҳ��g�A�����Ɗ�S��Tc%�C0��π��8ިht���6��-]+H��~�<>�'���eA�X�jᛇ�S�ڛ'.�@\��������֏��
t�ܣ>ߠ��tnD��8���Ӄo����f^��K�ݲ����
m��F��vy����<��>I��z���1c��v���>�r] :�|������I�G>f��	�?f~Bp�(�=�>�����ʛ\�ܟ���h��9#)���屙���8�@�+�����/��bח
엲y�W,�B����%z,�������=)��Y���Σ���-�l�v�{eA"Y~� ��e�_X�u��+�l����ֽg+�xc\��cn.h̳�����\z� A�X�h�ƿH}$�_���7���A"6=wF�T/Z{�l���.9��R��'�tfz����.6��!�з���g���ͺ7�y���k�7���x�N���%�Il��7��˧c@��0���<���m�C_�Л�<��FA�*t�V���������Í�O��v���ɂL�̹�qS(�������6l1]��^��P��y}z���������)��_U=fȍ=�Ytz�jX�Н��)}��󸴱����.�wpbKb:���YyXA1%�]�ą�`�͈ew�t8B#J
�w�%TĖ�&��i���5õ�F:������g�v�?�@6�>bk��u#��d�`4U@2%:��3g�GX[Z�kz�%L*�A��z���J��@�g�S����>�kڧ�onv���au(FˈY<���٩�J����(9�������ߢ�>�ԭAh���L�M����C=N��~�>���B_��C����x3�Ӡ��u�'��Ct;�>��Y��-֔>(+++�74����6t��/�$r]n�(e�vz��pŧ		�|��Al��^��4Md�1��>�c�@bK�R<�^UʑLW^af���s,�΀!-�mp@偼r��i���ag��N��X�r$�[&ۈ���!rlESW@�����I�,d�r\IO~Kk�^� �C�6&�7�d�"�j�^Sv}�T�C�U�rDFo607@�^7�Q8���%ZwF���v��ve�6T�]��P4�&b��=6^o�1aӕ��N�TSH�7ȍ�K���C�G߈�C��?l���S��p�� ��:[�0iK���{7\��MW(B�yG4�w�f�*t���H��m��vъ��^ ���2dVCe�
��F�$��n9Ah�$����M�F6$��I	�9PQ�5�1���@V'��et�M��O�������ꁇwp�hPup��M�1HД�Ԋ�- ��q��UBr�Uf�}v� @jg��}�#�G{{$���z����%��Ӳ�q4�n�۸�0�%��o����
�0W>xZ�Lвd�G>=J؀+x<��[�Լ1�3&!��bz�D��*��O=yKqH���(ܮ?����B�
Fv5!b�C7&���v���^N"V�թ�����R�>�Vԁ�F7-L�+v�oY�x�3�[ b�G��� ��`L��:o�ʽ;h�愞[d/��د2?I
�t)��E�b^h8�`����Tm%<U�I�B�u^Feӕ��#@$ ��t�VI5{��ʢ���v*Q�=^"��?0��-߭�3��kd���0W샷�!�y��TE�n�BI[�q���{x1�����Z��K]q������kz��	\ۂޚ�ϷF."ý�����F
ĥ���gF_H5:� ]��h`s5���)��E���M���i^G
-�KC�u��Vg��j\���W
gZ��j���z�����Zc�Ak,C��x�o�g��(���_��o|���?�� C�~ߦ��~�_��z��F���'��P�Y/�;^{�έ�wgź�u0�����}�'F̆�d`n�`|�¤�,NYna?�U��^�G�]����~���ZE�U9c�A��{�Q�U�X�jM+���|W��8�&��P5�~__�^^��+���m���y�y(L�]jP��#�m�5b��%I�Q�,�yk���1Sbd�>��
k%DsbP�2��hMEڨ��Ʀ8"E��?�n֕@y����^3�8����sah�ۥU4C�	m#�]x���H�ڽ�j�NƏ���6lWl_>�9KK{Q<��Z��|f�-!�M���P�~�9N'��Z�h���Bm}Y�U����q�)�Iw���
���pUk(OL�Z��}8��q���>��9��R��q���\�g���*7�z�l_rہx��5�z�,z�P(d
�B�Xzɲ����=��}�kq�yaP�
nL[BF�R�K�oI�)^���Z�M��C-���}��t�4S���5J2O�%Q��;����C��k��iB�ˈ��Wi0���J�y~~D�?��%F���@=K��i�#���`k�^��_y�
�)�au8-zzY� �0w�������Ծ���>>��b�(���S�-y�I� ��2��]+�G��Zc����D$�"��i��u�l�w4����
^kT�	�*�J������iIM֏��Q��ݜá�i�m�[�$EL��i����U���O!�oI:��}�]�7��Ơ�����K��4~�i;%�q�^����=��/!�f�dt4�C)%�s��+]���y_����b�H+�����y#&ed�Q4��S1-���1a�}YrG'��MmD,�[wv~�}R�8W�I�g=')���D����V���[�?�������=�L���T�-���q�::�"�?S��n�r�4y��x��<`?Y�M�}��)�FVlӌ~M-,��B�Ѭ�0R	E-̜S���
�K���*͵�V�)�(��>C��;H���9{�L��g�φr�SC@4�C���t�F�����PK�(k����˭�קvܜ'�˼����!���jS������oDbP��''�	�/��Ͻb�LEH�S
!�L�]�?Z�eH��01�f��u�� ���mFLz� ނ"�v>�je��.��o�L�{ќ3&J��k6�s����D�G�K&���n.��&X�O��K&SJ�����B�� ���n���Ϧ�����q ����n�ԣWŋ����ss�S�d��ŐѼ{W��`�Q_N�D�R��H��WZm��?^�t�6ӕ3A������������G��T3a���ђ{��\�ۤ��񺤐|�����`ɿ���g�R!Ww�2�����>�lJwg�7�q3@�����>M,�?��F�R�G�/���.FɏY2]�go��
M`���,���k�Qg���sww�P�!�u����؅z�2�%Lr�4 Ӻd^��<�q���ǚt�?�
�h	1���F�u�����Xn���4�l����B��8�i�4Ł��ꡯ-�R|�ǯ���+�]S���n̜e&��
���.���dH�t�۽ܿ@�$�HW(^}��e�dm��5L+�!�X�?H��.��0ҋ��	V���<_��*[J��m���3`14@k� �!�	���GH�N��0XK&����M'��P�%����@]�_RP����2�#81..�.I1�P�H��1Pt����I�R9��]�����e�t:]�Ju���͘����S��(�U�#�����@!�5[[��\��e��V�V\%.���+����_��!���^�?�K�=�b�~�;}v��^�"��Bo�P2��`��AH+���X<r����L�5����F��a�����!��ZG��RD�m���H�k����6��l��J8�P�]
�xM��Hֻe1Y�g�A���܊������AҐ2F��E[T�ŊTA������o���P5�I+����d�M��Hf&
�s,K��	�s�W���:7v�}Gq�@U"XUh@�ǋ�?}����L�5��RA���g��éB�i��Z� �(J}�R$|�j�}%�|��!�ƣA���Q��C�������/��@��p��ao=y/s��8�9��9�y�RHBD���fE�Gx���ѡњpg*��M��un��f����-�"���g���aC���a/����,N�*�
���z(,_��JY���s��a���ʘ��$'-���sK���1���g���Li��n1#p�:l
I��H�ۻ\����<��LusC3$�	a��u��.h��/yo����Ý��B�	�b��r����`�ʍvY_꾆�'����4u���]]H�¶a�	r��傿=Is
���-�^�lt������=�~��V�k!�	�gm!��W�W��\��'���I��@x�����|}�׀�kh-�u�V\�'>�o� ߝS)�^B_�V{�)�^��{�0n�x#��{�oV��u���Р���c�c���VA�A���O�`���ڪˋf�V��-�I�a9l�^�x�[S��Ln-�9N:����XdQ�������c$���ĝ���H	'�59AͤS�B�%�TX����(�5Eu�\��{<C72R�-�q��t��PЁ�Ӿ���5߯�&�b�A\�qm�9�oֱ�B�����c�y"䉐'B�y"䉐'B��}�լ����P�����'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"��OF^��@p��ۇ���y���!e����'UL�t��=�#�<S�/�]���l�૎��f{�g��?
m���E[1�;zVγ2ӠfȔ[7s�o?lj،�g
|}K���&ZVUӧ'5S����?^9A������W�b3��
�"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"���������H/��"���P�<�Dȃ����
�3�M��M�0���+[5=H,o2�l�Ӭ�ikuo��j�l�9Pζ�O�huX���i�i��Р�x�a����Q�)��&h>�Ѝ�\�>?m+���|m�&�o~� L<P[J�'�s����N�QۧfC��/C�_�6YP\�:K�Ng���`gY!V�?|p���� �Jx_�}0L�s��v�7B#_6޻��Ζi�M��
��&�	����E�I:IPpߍ8$֟8$)�ȫ!O�<�D�!O�<�D�!O�<�D�!���@L�d�yR��B�C�P�i ��VJث/��d���\�\>��ݶ�w��A'aC�l�����І�����3�'?��v3Wa���{VH�?�%,[j!U8\\gB�(�X��;B80U2���坙���(��d<_�<���#�eÿBGzD(�Pd�D�!O�<�D�!O�<�D�!O�<�D�!O�<�D�!O�<�D�!O�<�D�!O�<���#�ݜЧ#� "�P��l�����طJ���7̲}����2�EQ;���{�&I�,=�ٲ,� Y��O���/%̞��H��v`fOa��	)���՞��w���{��o����;7�j/�dYdn����ˮpf�b�El�o�Yq��|R�6b��~�
6y��Ź��'B�B�	yJ��D�!O�<�D�!O�<�D�!O�<�D�!O�<��o!o�eN�)��:/�`�?��.J������l�ߖJ�BP?�?��sj��YST���y���,o>�.�5����&�Q�4�g��Ds_sE;5!�l;t�[�F!O�<�D�!��*m=�_� B��"�'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐'B�y"䉐���;����m�b�*�V�ZpjTd�u�VTp D�`U��
2C""`EE�(�8� DE@��
Jd�L�����G�-~��}ﾮ�M'k?{�{��	tttttޗ8�VI������O�=G|I�����c٤��*U���#��a���7�Vǳ�/���5��d��JK�u���ڎ�ooN�&�f�ݿ���*���O���y�&�P��+ݓ}�}�8�j�t��-�_鼛�'~� ���?�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<���λ��Px� ���?�<�<�<�<��e��#e����Ǐ(Ժ}�a���Mfy��������u�;u�h<�r���E���k~�S�?�];�1�p����>�_�GN!Řr����Vv_�ґ�ih��[��3^B�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A�A��<|v��^ �B�B����������������������������������c������c��mŶp���V�|�s��9zfX�����3�+�lg��<��_�����I\���W�Y��v	��}���=��B�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<��/��Op�Xxak�b`���")�ٟ�����$�t����&2+����̟$�=f��3[�Z�.�������I{�n��
{��͔��@$|���m�Lo������?�h���y��֏���y��+�M���� 4�}����`d �RϺ�������Ü�t�����os&|��������3݆9��*�?Y~7���TI�7�o��_���{l[�n޳�QI��_�)�?��3�[+tč�\ �E�E�������������������������������������������)_�H��]��"�~���S#�q�ͣw�+N�2���z���[ߥ�Jw�����4.�@,#���ap]��μ~Ƹkl˟ܣ#&RcQD¾|5���u���?��?3nWVVv��|\��~�Ҋ:l��$�7Qj�_wJ{��+�.q9�#�A�u��W�����'p�]^,2ӱ�]9ayd�(��T5�ݐ/Ndy=e̓���<�������ɤ�p��ٟ�#
7�=��}��H��/�<(!�~@̷��r������Ԛ�Z훬UK��9I����\P�ݵ��r��'���"K����iS_�a���V_l뇱����؟���AoeWv���:�R��>�%_���0����&���u.4HV�Rg�hS�;��Ü:�9H-��iZ��ۡ�3v��e�b^j�ӭ�$�444��tn��0'����8e�C6�g�P�����.���:��BK�-�i#�K�]Tfk�m�7Icޞ���Cq!�Rd8�s��^��dr _ˁ�f�
Ě;Ŋ{7�<f����D�u�|��?6��k�Xo���>߀� ��q��+�L��<��Xa���8b�0s�XtV�(O�_��ȋ�D�������1��k�v�(�7F����8̠
$�7Gw�IHۍ}9�j��!���d�K�ܥ��v��-��������o�Y��L9��̾=��:L.P�R���eG	��I�n5������"�>���j�d�O��{�S ���چ����O�b�=3��yQ�Á��!֥)i,we���,{[J�bK\�$�Uν����U">����Y�;�)���2�����V̳c�m�2���=�W�X10 �~���l\9��d����Ք��M�K��_z���F,w	��X-Z���~븸��O9����(SIԴr��Ĕ�O���{��Y��HV[�~|��3�N��r8�� 'ҧ��׍Gb;y��/��:1��?vx;������dIu+�O���h�T�7�2���&�a�tǿ;S}ƼO'6� �5m�������W���jZ��P�BI$��{�o�c@��xv�5v��5ꙇ7q[:����+1�Y���� ?��モ.�� y������!�<��i{e�z�O�H�#%�]v���?rq.��N�z:���ð��η0aس��M&0�����x�x8�}�[�I��ڭH��.���@!/���O�����1�%]ϭ�kN�mi�yź~2�F�gq����rQ_�߁���5�F딬���#��_#���נ �k�t!����v�2;'�3Tt�Uc��ᶅ>Y�& �7����^ ���E�$8K(��R����X�~����\���w7�qOV�N��ǳ������w�c6q����}�ߕ̰1���OBA�|$�em��ԧ�f�����\�A(
�@�8k�J�쨅Kh�RFO4��%~�K��U҃���ӭ��bW�}nV�=>�&8^�	L�7b���e/�0s��_� �����N��Z�Ip�+���3~K�V�*LG6�R��z�?"�a��,�@Q��at�2G�˿������`���<�����o��sO�����GN�:���ot�1�{���#��ާ�����U;����cY��Q{th#�ژI1ɶ�#>��`��I���C��%ˑS�x��'>ܮݿ)l����C~�uv���p-â�灘Y~�?�"6jq}&7���:LN|����*�/���pa�Wb�$�5w(�ܶGN�O੾.�ᶼ�M�u|oyo����@PV�CNbf�Y�#��=��o�E̬�g+0 7�ߛ���O�pE�J���9��F��+�S�x��)�x�2y���ȯ�?ڵv���AS
��q0��Y���M=hr�p��[��f<�|cfЎG�Ev����_gL�gR5��R&��Z���*:�gDjk�*�\3�uG�,�
����?C�3����a��N�dY�T#7l���oO/�P�q�(er"f��ȯ�K���C��C�� f�@Ѐ��(�����A7��A�@��J h��J h�����w��i/b컽 Cb�C��A�@	��@�@	��@�@��n�7��A�@��J h��J h����A�@��*n4Pq���(���(���.l4Pq����T� h��J h��J&��&�̯�@g��� �)L�0��d�.�®%�kC�vm����7(���(�����A7��A�@��J h��J h����A�@��*n4Pq���(�����E����l�<)k���-�۞��Udn>��A3k��f�d��-���ZudN`�U<�uT?�~���2pt9�磕H$��Iq���)�����#[g�֡��<��@��?�eހDt�OF���v�y��n/��P����\�^]��F�ޜ*���O�<�q�x>�7r��:�8Zn��]�����bG��s���?�hl{1���_�o�~0u��y��x�(>j����΂�#Z�xL���N�O�W)�aփ�j�ȼ:�C^�5x�΁�]�yDKT���B����?X�ґy��C^�=x���D�����
q�W��\�`��G�Րy3z����u���V���^�ܡ�u:��:ޏ�t|Ѩ@�@	�@�@	�@�@g�iA5*4P�A%4PA%4PA�	 h��!Ԩ@�@�
�@�@	�@�@	t&������K2��w|Qy�Ё(�Ё(�Ё(�Ё�����J�@�@	�@�@	�@�@	�C�@8�@�@	�@�@	�@�@	�C�@8�@�@	�@�@	�@�@�h���������A�@OI�Q�Ё(�Ё(�Ё��+�1*��7@c���I�j�	�&���j��?�&�mE	l[Q�V�|M�����M��5��UUc����S%�����Ǿz�|E�U}�{ ���ˬS j-���RG\���9�OBB�W����X�/�L�<TZ���Z`0[���W��h�]��"@�1unGFi�H JHoX����ٖ,��q)����݊�	£,?��QIvO��W?o~��~N����>CX �,H�����T��H��y3�FD��ɾ�V��'JK*N�q��w�ʸ O��8��VPI#b��8Q`
2�ܗ f>V��(ͩ@%oa�~�tۻ|�d3���g�Gbb����9*�2�(���9+ q��_�e���5�*e��\���QJ�40�ho2�C��.>����;TSG��
�Y��w�ʸ ��N�t�*xT��*q*HWJ�ϊ
�y.Ayt�`:A��74�<bc��r嚝�'�0��Ғ ����Q�Y�nOtvAFhx|_)�OeW!IE��c��Q��8���޴��G�4/�c�bɝ{ٙ����[>��Q��/�(x��ۧ�8_���4"^h!���:���V�pI�����r�|0Q#��L��:�`(��稌�0�j9��� ;�F�w�����abh�'S��RQ�~>���_b~6 l�h���~�W����_������A�!x��Z x���%<�ц��h����6��@�@�t�!l��:�6Pa-6�ц��h����6��@�@G�J l��:�6Pa-6�ц���h���&���^�_	�]� x��Z x��Z x����ׁǈa]� l��Z l��Z l�K��@�@�tQ���h���h���.U6Pa-6�E�J l��J l���T�l�����n/��#��C�@	�@�@G�J x��:�<D���T���f�S��	a}�T��e?Ͼ����o����w�m��xg������C��f��;������&|�hՆ>p���$�
N�M���F�3j���}Z��������z�Yx�9�kB:���5r�͜h�M�}6 ��V�'��=6ra�qe������@3���݃GN��)�M�����G���D��]�y��9�;:�4�y��W@3���Ǵ�>�dC�)�I��TG�����g�?���5kF<K�P�5�,b�juGN��? y��Y��h�_+��v�ܗmk��9�<A\�k�f�9����v�S~��=C@5c��o��Q�̃�'M&ǹ/�r}T{�+����/w�|��3�����8 ����W��a���6�\M�jdMW���k�u�a؊#wt�ȢA�x'6�	�J l��:�@�@	�t����h���N06Pa-6�	�J�{`#���5��@��hC�@	t��<&��RK�u����WX^ay��
�z����` l��:�@�@	��@�@'(����a%6�	�J l��:�@�@	��@�@'(� ��I���/���>0�@�@�!x��Z x��<>)6����h���>0��@�@��@�@��!l��Z l�a%6�a%6�a}`(������ �v�
\5I��,�;�M�Ki۔�<r�75cq�K�
_�0����V��w�o�3��(y� ����#z'xGg �*I����v��ޑ~㝁g��F�;�{��ȏ�wމF�l��#i0��_�a�>_ ��@�� �����*��b�;L5�����w{��u.2�p_���_ ��7�z���т�(huZ� Z#��8A�������/�V�7�:���т�����b���I�y\�$\ޣZ	���_���z_ �VЪ? ��U�������=���{��a���W�j_����U����@+}��5�=���ZY Z��;	?%���_�[6x_ �~�:} Z�FZ��Ck���Z->�n?��	��~ �3�޷l@����A���6���6��@�@��� l���D6Pa-6�&���h���6��@�@��J l���D6Pa-6�&�����a��j!�n/ ��-<P�-<�I�J x��r��4��@�@��@�@˗�Ʊ,G6�0k���lQP[��-�EA'iآ��Z l��Z l��4��@�@�t������l�O��w{>�_<��}`(���>0�!x��������@�@��!l����6�����C�@	����dޮ?cR�t��2ww>���i����Ic~�t���o�̾�?v�W�2߮���D�Ȥ��0Qc�{wDG^�,�kR�a��0-�I]��̜���!t��]� �%+�No����:�AJ�����~�W��WH���O�Ŷ�X�+��bԋ�>��t\VR��\�F�O[-/��7Zi�x�i+/#�|Ƥ�jv���%�0&0&0&0&0&0&0&0&0&0&0&0&_'&G.���^ ����1!�YU<�����M-���"�Ŷ"o��kO.fdw���'��i8bx�%�R@@@���G�5�8$��u��#o����9t��d��47��ȭ��Y�痦|����8uu�ӊ>݅�S��⻙X�f���M�Nn������WT����:�"F�RV�G�Q��>7�fi�J#u5>OP�<�%�g�,�e��b��r�����0����g�|b�;e��r\S`�f���~A��&wK$T�{8k�0��'P�W���g�u�nM���i����arzb��>�����.N<�=P��g��� ��4��\#rz)���Oz�St����d�,=�2����':}��+8�t	=}�a��(;��m��緊D[3-�=յ}���d�e>�����I�Y�t!Y(��cf����ҹj8��]��ˎ���bM�������d��C�u9푴֬�/� �녙%C�ͱ�#��{�J���������b'�w�U3Xv��i�j{$X���T�!��B��A����?����T���t�e�c��H�׿yv�0+����U��k!&nV��V��H�x0�	��>f�4%�������)��D�����\�d���g���|�MTҫ��ӻ��FQ��W�X�gO�R���=�˓\��+�P�!�Ņ�vQK�f�;��^�Z�sXJ$�Г��5���j�55BA/{c�~B���{/�CO�e�}��a3'軴��w��_gzY�)׊47G��!E��YEw�V*߳�<ƴSriE�#�.���~juŶ��'G��o�7ǧ�9�a��Ө	����-]\x͠�t^��#r(F�v�W�J����)�����w����7���G�
���q!�?��ECr�0n���6+U��g�]>̕�&��GdG�.��Ѭ\���+g��'X'��-�.�lˡZ����t76���FtR�֨�唌����٨��&��I������+����[Jz��;�E|&v��igΊ���K��

������	9i��s@���	��H�B�TT�Ǐ���G�G`J�WSõC@
�|�d���*���ҪXQ��z+�-U��f�fD�Q**Ǔv�	�d�S��	��p�u%�Rs�}uji~�+�ֲŭ�g]�"{�=�S���L������H���9��$�5t?�bt���?��h���/,�j��^���,~E^��?+����^��d[l���@&��� ��R��e��n�C����}�����_��iL�"58t���%m����t]� k��rI�t۷e�ж湪�rN`��Y�z��F.y�-G�J-�i;r2v�m�:�sm-����l�W��Z�x��<���tZ�5˴`\��W�.���Q�N�BV�M�f�؇:���sA�*F릎�R�a�M����{�/ܡ~�hV�h�Y�I�'��T��+���� #��ۧ,teD��u]%��!��<Ž��֔���a,<�����k�%�}�`r"D����@nr����7��jf��sQt$�R��U������&�]lI��W���62K�=.i�Y!	��?ϓ�K:Μj���+8ĵ5N#n-=�3X�̌��	N2��T�G�#]�r1}�:B,=�#�gU�����I��;��G�{q�mS5�sO)�v{��m�������{�5�q?-��n�H�����3믐�;iˁ�ʊon0��[�뵆�����A�=�1}7r����p;�<��-���Sn����VJL��I]� F���4�n&��߬A���p��h��۞�����v�\D�u��[[]'���+�v�S��hyݐ��������A2hn�'֡�s�NɳSG�b�6�.��p�)iGr<Y����Q-�g�p~<$Fj����3p>=�f��k���jC��(v�Z���T��j�u\�����ԅ�G�f4.RPq\����㰘s��g�xqF-1(CuHU^�(7XJ�J3��i�¯&C��r��w���Y�Ⓗ����PT�(!�xg�`�A7&�b�7+��E���Ẹ&�(#l��̉8���ͰC��&Rq&���0Q�y̪���L���:���Ɲh��V��7p=��&��"Ucy�uwNmO�H�\0�1�ڀ� ��5G��ew�)E<#l@�74jy_��ޚ�w��8�>��<�$X���_И��h�O�s�y��&�z�C��3I�5�:�zj�:�;&d�
��V��8Qa<��|r�$�қHj8��sL�Կ��~;�uK�\�ۉ�.F��`��� �p�8���B��ӫ_=k}%�h�:�e28y>��qP
��X;R�1^�'@������ ?���ݹ�n�u1�t-���C Oۼ�=N<w)$N4:�+�dx�Íd/�ޗ�������0{ͺ'�sj�5@�蹕�[#�M.�֚���%P�N�aֵ�ۻ�g�3�Oi��%�@Hd�*⦍�$E>9ڬ��e�3~^Ƣ�0�
\E��3;�Km�����c�9���Y�Ue�=�DB��t��-�
Һ��\�j[`�j`!��?h���0̦�o��:�znױN&ە��ZO)h����ʦJ���ls&�w�~I������a~�p���v?�,�o�8�ikB����#y��~��4���'���æ!��=6� omE´n\��`ݲ�P=N�3�V7�e����0#���d���\E*�4��s]�]�}��[@%�[�9��%�a��}bO�i�I3�O���������+v]*l5/��:��K�on�H��v~W�#���m݆���ٯ�9�	�{�����O����鑛Aw��G�7b���7b;+^o�9��4��3W�8եu]������ �V�=�JW���_�a<..գ�i����f��ka���[
��bC
�-���i�}��Ϋ��n	:��xE7I�Lf����g�^��ލ\��m ���-qU�R�i	�;S�D�����Aj��+*���\�=[�f����c1���i��n�斊�d��3N>ʘYj�|݊-.����85�a�oO+-y�L�K���-2�a���U��G�X���Ӿ���87��,k��[&c.�\֡�`�5q�C 5��}��!p	�tp��U͐�rRDO�+����%NO���q!"H�m�_B�|B.?��O;��I%<��5��qm��n,:�kurڶP���׃LI���s����G�(���H�eV�5�k�������>��m�qQ�2�FU���W�0;������M��%HUa�[�o[jd�s�Z��ObJ6�Y��������c3��'���y����.7AG�CF ݡ���gK!N�����,~��/H��eGK����>  ΥW��T�������bGuw����є�'����(f{�vϞ�>�3g�\� �����] *�@]�m�:�O���v�;vp}Ϫq ^��h�̂!�� y�'�Aлd�/��#�#S�p ?פ��̱x�7O��zsA��l�s$Q����r�dBwSa�����^n��-����ܜ�2�g?�'�ީiH�hm�#$� V�ަ�b�:i��� ��`��Ԑ׆�1E9�:��夼�ud��?*l� ��mb�x}j����҉���&kWu2������+�/6���.����q����F�O�xy���5H
Y6�1�����^�#��"ܾu��R��v�� ֥�G_?�P��Y�i���NI�5oY��r\m��$;s��C�O���g�D��V3K�ykM;o\Y{�� \���4����U����ry�� �rg���(��_y�Z��$���X�(vK 
/���r�M�ƣ��3��C+&y����_A�k����{#)��|Z��.�X���raѐ>P�x���T_�῿��pΟv��YMY/��-��ui��6�n-��r���Z�.0�����~�
��[��*NX�_�����z�J�c����s�^��V֡	=�߲�ϑ�#�:Rش�Օ�h�Z�x����]Z@�f0%�ZD�wŽ���+����uFuU�q�E~nNk$&&�h���I���N�Ύ�{H/�=��r�*�}�g�I?�_1�T'��c�9^M!j���|�R���ݦR�\���+w��H�~+>]%���m�|1��� ^z�%r3�����2@_�u��/6v:��Y����bdgc���T�������~�	gR�_�λJ�/.I�Ǟ���?K�R)�qN?`��Q'륂�L�R��
L��r*墴NLr$K�k����9>�Bj�H�cg��� O��Gk�s:����/�����7V�\ J7��z7ȸL\`�L�گ���^���Q{K�Z3���Nn�n.n�����Ӻ��ڲ��|F���Z��}&=Y9q;��'��bob��L���ֳ8(ܞhcbV�0��(�2�֌�"�\���:�Y�5=��:�!%b�
�o'b� ]��D���m6v��:�`Gr����r����m�	��]@ӌ䎼@c�Ãs}@��9��et5�-FV�2�j���"W+�Y��^#Xj�����Y�C��{~���õ5t�^�m����ի��7ED�rn\?cƌugL�OMS�9]/:5�g�	 *�|�U�E�>9l�U�\ԛ����K��9G��N-4\�99�tl�K���A���Z HB(!�Ӽ�@����'V���2�YF��L<�F���D;�L���K:7�j�`��&�u�L�v���x�O�`��RM���TF���BA�ȝkp�h���j���c�%YK��F�MDޮ��2MK g̘>�)�E��K�:�� ��5Z���X�r'P�V�7ؑ`�������_ן�*��U�!Yn7贩�|��d?_d����Ei�
���^C��9ǻsdq�7��Vk5��\�� �y���TI�3\��֒���R�J��'�ַ;��۝�:#����:u�i.�ל���g�ą�i�"��M4/�������IDAl�?֌tS�}o�.�[+R5��O�8q}�ᅣ8|�*�@�Hjp�+ O��-#t���8~��(�J#Eo4��G!����I���#����Z��}u�E����N&�!?$yu]�A�|Z��EJR݄�թ�{�Xߝ{��CJ~����������������o'ά����i.]zN 扬�P���mi�a!�\�t�~�ط�%��Ճ�6��6��]���Sś��U��=��`��rP]�$w`�qaj��t E�����:<s���6C�"�4B�ꬑV����G-��6p#�D���D�P��f�,:H��'z-�F2Ťd/����xαe���J���2�:m��S����[�W1r#6T��q�t����dKc�s�u��Nf��VF8���޲%�4O�`a�Qpu�c�>�@�S{`=�F���3<�3y,Jd��ȯW�&�Op���y���]���Τ��Y�s7@ڞ��1q�^dT����������in�r()�f�MJqx[p~Z�]�n��lbc�I�
�s%-�`���2.ū�vt���Y|sC�,�ƭ�/��� ���An�v���T��þ�kn�P��-&mͅ��q����u�ֲ�r��i㉬�ߒ��J�s7�tH��5�����#�U�s�b�e �;r.�4~�ah�6F���Ĭ����΀�����>����ͳ<�`E _$~��Dv����C�ұ@�df�/k�n�r3��;X�f�����"o�p���;�~���D��홧6~�$| ��R���f09��A�T�Y�W4�M"���%��=j�ߐ^�R�G�յAZ�̓��u1���� �����9�-��bA|)�	���Si�O�Sp;�+�b=#��nxf�~�>�8׎s$�,�t�ٟ6��U�,�����0^�[s��лY�񏏚�o��0�d"&x������J=�o���T>�y�6����}�t�h6�є�N��n0O�Tqa-?x� ��l)J�~�����Ձ�zl@,����~�s�7��Z�-������X�橤��|��-�4⹄jl�j�]�=��G�`\'����iГ�!����*;�@�k"��}��HM矺S�fєe��ci�1Q쵤�)K�h��X<p�D�Lx;��	�-�jm2Qm��W�qWo�Z��{�4��,��Eꅻ�����3v�G�}@���� "�_|��8�Vb�9R���T���vF6�������b�XG�q�V�lf��@D#Z�("K��ŭR� � 
/"�"��U����)����j~rR������ȀOE���6����쳘 ��^I;�!tf0+m�I���j��_.}�1��,�y��jF��!L��BZi3���C�(a��Y�/��D�M���Jm�
�@SP�Ʃ�bE�y���	���E�W�c��h��4�ͿP�� iq܎���ul��������1$v=טBP��� j�@+��f��fɯ,���S��=o	r�c�F����7�[q����j�ܮ69͹�YR&���*H�xl�,�Ca�-9��zoN���&\���`J�k�[-�X��%o.�i����߱IB��:T���o� �N�\�;X�B����N�̤dp2!i�w�Mv�J�UW?� �������ԏ�j�%�sA�t�|�t-��q��.��� �W%�@��X �a.�ܻ=�t'-�˸��_��b���.��/A=����H��6�x�Q��Ky�YӸ���V�Gf�֦�V���fƴ��%1�[���s�U�1药NL�l��n�i����ۓ��ض��H =ymI�3��b�*��=���6(hTt��f �^y&�t;��5R��&�Ӑe������g�eu�g=l\�aAjs�Y#���]�t�{
d۽tO��;���OLw�-�]��Y�-9�Q��=��-W��ޙY׮�����b �	fx_ѢoR�}�7�WD]��ǚ�`�uT=}��l��z;%�-���=t�2�ׯzCƸ\�e�(9D��/��ܟU�O��A.��֔��-l�K�ŉo;zà����f�䔚��ws��d��,:
6�L�W�Nu���s�A+��Ð��?��ӽ��D[T��իW���XR� #�7��0�\���!�,����b�Dn�;w��r��g�n,�5����,�8b����\˻+�i��hDȪ�fH��@E�Ż������<^�ɳX�������ݚ�fG��q��b�e2&��j
n�`�.�����.5
��a�Cof���C͛��T-���f�dh�b�F�:2o���2fk�,�'�i7��m��|
�֎6L��*&wmдa&�)�ɋe��a.�-v}���ӫ�+Xښ�x�z������̮%Q��D�2��^����2[Jc��m��#b|��ƚm�_��M��⁙�vJM���z}�ӯ�E��/kD/�v���!�=��ޗTY"[��;�vJ	���7hƘ�.�����O��Q������pQ�}����`E��17!._�[�S�n;i|��@�Ip�Z�%=��4�F�P���0��KmJKU��l�cO32:���@�_^)�H�{.���9�0�㵜L2����ȿn��2A!U�?J0�-N�UK�*6��e���>`^��@'4�Y}�D���o�ؑ���BaŁY�5Q���|K$\��Po���#j���A怢���
�,���<zo�KiQ$��SYkWV�=��E����n|~��WB����&���Ɔ8�-�q���n3;Bg���ړ<X{8U-����;��s��TR�8�`��}�><�<��5i7��������V]w��士� ��ýe�`�=��w" ͒�E[��=�R�c=��'k���-]^�u��؈����n	�vs��s|[ܱ&�XGk�u�) ]��i|AG����<l��oxH�/�: Y����Se�O1���	���9����x.���^�Z�ٴS�x�	Yk];o��Vn]�~�)�M��7)Z=�T�q>=&<��i�;%cL{v �F�%w`�=AL��0��3��~K�Y�Ys�%�p�9�v���~d��N-�I,B��|ʖH�~\0���%�'>#�I���	����zw9t/�K�Tۤ��P��f�;�rD� )���倇�Ǿ�܀GB1�����kq۔��:(��:�qS.G"���'��y>P�	�S;־�=�����cF��M�w�Z3�+��@8=@8ש����|�Y츐��U�l��m=�5B��S)��i���wn~s+�P3v�h���,ˑ�결�%���1�@�{Z�����ŝ�k��9O��-������xa����ct�#����D0�,�3zzhCb#P)����}ϣ���\�r.{�'�m���`yi �%���z܈2����	5�.�xu�;���$�~�z{�t�k�v�����(vGqC��҅Q���
yKH8ޜʘ�O�1�٣�9��q1�!?$�̙3v����m�	�d���P�2�H�>b�'��T�^��x���x�tb��0�����Lw���,�)�G�����":ӬY�A��0��խ&��J��㜩�rB=A��p�/|�v��I{ݶ[]�vq��5���&�˝?c�����{N嗀�2�jk���K�7�J$&��ky�I��K;s�@�B��t4�E'k�M#,֬��UZk���b@}�X��=�g��zPH7�0#�=�A¸1�L��ST���;��cS��GW���T�V��4ߎ)q��FA(R\6��^D���K��~�'��n���b u��~z�J�w6�Np��\���r�v�.dd�7��oaU��ݛ���`2t(d��,=�S����+�Q�$�6j�;�UbN�kT�dLJ����.6
��d�~���{R���J2{����/܁vU�f���
�җ �x�z�]�������]�p>�JRZڭ�$A���ձUMy&Aąf�� �e�C��O��mi��2�[bțؾ[��z/<7��`�GcӉI�)�l�J�X�e&.q�ܹ���������q�������5�y2���S�M������0�U���|3�뼅��V�a. ɰ)�in�e���.j����f��}T;Ҝ$��S�R)n�3��o�P��S�z۞.I�s=j6��i�'�(��������.4���5���t\��"(y\��/��:�a:NH�g>AVU����`�Z�>���i�)dM���ć岳7#Y>w���W��=���X��I��EKu���J:��~	��rKH��F�8�xРmP�"rj���SZK�o>��ܶ�MXyq'�����Zp ��Gk�e�d"x��~�d�;�	?�^P���Bp~�n�w����XFj��d+a	T=�$vs|����z'x3�e7 �H/\�yYP߰�;��1��j$~j��V9�� )FD^��Ij�3��3��fd�h����D�a<ť�lQ��;�4�L{wi�ЖD�vc�M���=}�g���/��M�%��88��H�����"���`ݣ�Nߩ��M~���FS�[jiD.� ks�-S��ٟl&3F4�������>kͽy�\٫⑞샰����6;\k5S2PZ��U�Ȗ'��{��J_��E	Ȟ%3�% ��מ��4�����ڷK�K�Vf����Y~��6^Z:��%At�jAY-�f�F��5#xJ!�`x���ġ����d$]���+��*3������}�^�vZD!�h�8��2j+荭c�H ��̩�y��i}�[��|.�����)��D��0��hK�P�t�������m�u,#\���6�u/�M�{��I����]��������A�
�~ �T��Rr��G ��BkZK��'��.n׼��������-��u����<�a�C�E��Zw���f��|�9��~�k����]��� <��ߐ0&C���7$4-����tͤ��в��	�+���g:-7'HV9]#�בV/t�x}.��U�k���#�K#���2��U�$��WLu��`��*������Q!7��>�nC%͓��}-X�R瞈�,�	٤��1X׶�G��d����Ϛ௔X�����j����j,�?|:t��0�\���?�U���h�o�#
\���a�eȕ��68L&Լ�M�f�C�:^���#��yPjA�YV�ۂM��q(�+�Km��q��'|^&Oy��!�q��s��)�2�N�~��,��A�-��
nEF�U�c�;��5j���bQ�U���r�֌��/���msB.C�0��i��?�E��9fSq{���3-�'�
*2|�r���J��E�rB#@�r�$����L�����ǫ��l��w�ҕ'^ϛXQ@�6���9T#j���:��*������b�`��s�O�������$:�Q�n�ǈ�/i1�k=�`��*ɀ�k���� G%P_!+D��%<k�%e��\���۟8d]ڃ�b��ҹX�z&r]�:�i�iO����k��]��z��3��p��I|4#S�F�)!����g�X�<�9�c�o%��_��eȵKϭ�G%!�>������5iW-���\/l��%��[��M�����E 4JWn�N�d@G��!fN�ϛ���U��A��R����������1.����q��LId�ڔ��CH�}"z`�n�`�l��o����v�1����7_p6>H�#�Ӑ���r.��L͢{�.`T͉e�:���#vB�������=�?�Wۀ��ﺖ�1��+Ȼ��~�ّ���`�p��6�9�����V�����e���.��g�gx�{����gR��(�xP\|�-�+���x�H���i*x�R%ݘ�	�~����m�l[�k���Ӗ�]�0=��ف�xM	d���	���d���H�g�A�ar��PPg^�-�����q�G��ӈ�pZ�#��xdo��G���@�O7i�������/���g�g�\�� h�gf���vf����ً����+�H=O��p>�*=���ˠ]���0�C�O*���T��
�,nG³�]VVV����Y��(��ґ��PO�,�c�\�o6�����ׇ���=|���s�xz����2��37"���d	�d��7��cF��*���0����ְ5�W�L��ΞBCns�^�(h��u)-��3ȑﯼ�Z�/4��)�+[�1�����*������Z3 � 0�N/lK��xG����g�(��˜";��N�Լ���,�_�3]��; !S�Ӓ�:M#���M���iu}�*��w$E�#�)*H�'�{��Q�����6���S�;�x�A�s���(u�ҥ�h i���>T��V��)�߂��4e~�tS���̺� ��ks���P]
��z�#��d+�����߯��R5R����5����H,��yo=K��ȯ:�;��\�iB3��Y���<��qC��PL6i�U��F�g���ĖR)���~�mJ�a%"�`Rd�{���:�����ᦣc��;�w��4��}��ϐ��mH����$��������l��J��v5Nݫ��Sϕ�]]��
;��!��9�N׀��5���^eG�H�`�ť�����d$�{耤�$};�т�er���>qt��q5���>q�:�x��n�3����A�*:-���Vj@��و<�"j5�v���c[��u˚EAΖ��/;fYT٪�|�^��p�r��=�io�9�Ò�L��a2� �׷A���<>u�f�V�@�}?q_p��e��6��m����Г�����ǫ3�bc��0���S�{��6�����ȭEv�>�������\P�t�������CI �g���
�Q�c��(os��J�(`V��	��m͘SQl���s�7:��{)�;l�K�@E�BEhN�]�E6G,ݺ��M��O�Y<|�����F�8dǝ���,�'�K-�����[	���!�wv�=�=H�z�	&B(�noe��������ǍiN癀dS�1�D� �M.���Q)�q���
Z27���~2��J�(�@{\,�9 ��=Z����&���(vO��$�S/�0�P����F�/������w�'�	�u9v4Q�.������T�R�͌ʧW�"�������@m�o��GfD�^Fn�k,�'�h�\�4�%LJJj����ՍEw*5��6Y�}��ꐄ�EI"�o��n�,S�K@u����q�U鎼��H��/)6]�ϑ�1P<Y��x��6���ǜ5P�YZ)��`c��O͘+{m@%���\ɠ�g��ǗĒA�����DR�뼇� M����[�����lv��G���r�?�m�������|��S�^��妻�K�ҭ$
�R0���C��xJ9.|����5��&�ke�2:m���qӸ)媖�+b&Ȫ�1�i��s�=-z��~S�h8}*i-�0FS�Ѝ�p��k�T�H�3Mz��u�Gi��e�a{�m��[�y���^�TfH]�������?x�sQ��y���\}?��t�N$���yy�g�V��-G��0pr�*������N4�Y7� �K	��8���TBu����"�X^���8����	m�4N:ys� ��Vz�WnK)��K"��4�C1�%;w��k���9�#K5��y��8�����!�[�1�:۔d�@8�R�:��8t;�ՙY�YJ���r�� ی�8]=�)��!4��7T��k��Iz�P�ac���e���nv�qs��!7���]o�Vt�H�\�yo�8���tI�:�GY���V/��役1���|���+������v��B��A7�!���"[P�@�K��O��r0Qݫ闼=�m[��Gޔ=�>�^<#5�,,�֯�J亍kYƎ�m��|O���k��8�i��B#:�k�K���J�B�Lu�J&��T��u(?�kq�:6n-��u�<�ٛnM��yP���e@�َ��,PB�{h8#���Do���Q^9Ї�Tؒ������k��ȃ��̏�!���Б<�ۙz��.]�g晄�3K����RL��5��'���#E|��>^U�3�vU[�MC�4 p^o�̞��;.f`��`�?��Y�!������9�������3s*f_D��{���;1%�B�[.}���b���A'�GWv�c[��MJ��̑}s���*SIqk-�뭩_K5�h�	�Y����O��ib�I��&1�:ڭ�Gq
r�s�^"Y,��s��K|��Ճ;>}���T�ک%p�&ҏ_��GSJ��[�N������\i��";H8G�$ާ�G�/3���:��*gtS�c��C#���'A�4E�J���sc۷c��-c�8��~��sd���I���zdۭmc�^�Af��G�&U��1|j������638/߲�͈�bV�"Բݱ,���M�D��]zZJ�߬��v�3x��M�Aa���l�bs�b��0�:���;s�����H�(;�\��$z��qԟ#�<�GP��.]�5��"��7@uK/w�Co�M[ϗ�h>"S��������X�O�ys�̙3�!���{�6a����yT�W��ZߢU�"Uq@���V��Q�I&!$)�����"��eH� � Dd���1@��9�
��Z{���?vu� �����~�>�<ۑ$�a��e���l>{����t8`��K_R��r�'2NO�� ^' �t��od�n{a�AD(����k�9�3��)����h_�Y�;�O�բ���������Ó@¼���z�]N��)�ug�$���ic�ܱ�"�-�YN�
�0�>�ӓV���E!<��"�I1�X�F�k[V�y��8S��P h|f�z��R*�0~�͞��R�($ � j#����N2������,�R�ǈ�o��j�P}��:�ͼ\Iz#�l�ڡW�|p�V�d7m Ҙo��H#/�@|a����H�O�e��VX� x��)����"�d��D�`�j���]dV��U+?ᡩ��nU�=�T�b��v���;v�NN굜'7�T�n�d4.Ƥ۞9����_Yl[a+֣Ŀg8��^�:�8�Ǹ������d��ш���~(�Y��f���;� ~v:�Q������	�g�������X�qvzNֻ���g{EU�Z�_k��|ƀJWw	@���sE�FT_���o�Q�@}(��e؍췬�W�9e���j#<:}��J���^w��
\��S�W�q�u�cƼ��35l�_�z���J�L��p�V���Bً�W����y��P{�a���C�eB�*���=!�<��kk~�?�^<���=[��s���Y"��i'.����=U.{^�I�o����@3q2�(m��D�G���H$OrWH��(��ZC��(5זk�&��D����0,=�Z��%��#���S!�B�0��绡9Ϊ�0�9-�yr�
 N~����.�N��O�:2����&�<�Q����S1����s�<L�о:F]j:�ELZI�,^@�h�'�j��4=\ؠ����^�~���{�
����6����n8:���O���*:��	�_p�4��t���S_6���z�:�pA$o&����)s�L�s���Y�IX��N�u�q.ER@�Z�G�AI��q�� �ث���.MW@d)��+c�ʻ<�<�|��Z�?��؏��DIrVC�T�Ff��~�ϧ4f;�z�c��|�K�kJRQx����U��?^Y�"�d�y���N�U�Oc'J�Kz�;YQ8�� $�Os�{g���֩�����	�c<S茰N����9�Bc�p���ĉO(\Pb���䴣�M���oR:(��ޠ��,���4�Y>���03���a���Jހ`U9�����ڬ��qZv�Z��J�諶$�6c��A�v-� K�]N��)�����Q�zx�4����J��T;�񀡝Ya�y|Ovq�h��0�|����o&Yv�?}*�r���R:2��u��.�ʋJ �����uUF���������7���$D@ÕW��Q\����=!������</�/v݅�5���2��ا�� �HL�_juO!p#lL9JQ��2	�%�|�ʨzi��L�N�a��]G�DNΤ6��q#�'�:���y?��z@:��+�zrW{4d��p3�o���O�uo�z�o���itx�Ҟ"3��N�x�cy�l_�<��t5�?(H��A�����P��
��_�gXC	���4x�����Ί��TB�ג�يS�'_ewBx�sz4�v���FA~�(��������?�;�^����.�$� ��+�N�{� �6�l�~M�f��d� ���P����|?!Ȁ�p4g'���ٕ�ߕ��|8ӎ���It�S�i�D�"k�v)˟<3��q]�Ͽ#�i,o2�o�a5�eI�L��q����
x;z"�{p>3Pp���V���lO�96�w�A��9z�3��]���څ���Y�Ѫ�ͩ��8Y̻y�/��*�a��u\0!+�6�n9��f�0��a�9�r��v��ͦ=���)�P�ԍ���=>|^�i�y͇?���t.�6��={���H�q���dhM�N�<6 �����.3��(��&3��@\<	6��AaU�z�K^u�L/)�E����B!��؈�E������q�'в녗w߅��bv9���!�͛��}�o\f�뫊/v��"�&��A>��d�-�U�&��#l뫎�tl/	l�~�Zs��b�����~P	�Eu�P���Mp�[(b 1��?����mO�_'�������ҏ�:��^�l0{���ū��o���NH�!����\&�����'r�
>�d#���`�ʍ�޳N$T�
πIݥ��(��ُ�oê�=�N%~ &}rA���x�H�Xg"(�
Ќ���u!6OB���D�C�,X$��N@�P@����H����Y>����/���H ��3r'軑���3�/���{�v�Y%)s�^ �i��WdE����Lu'Arr�/v�H�>�N�s�p挥�g����6�`k�<�ݤ�6��&^���Wd�M��n\�_���ZP/;�B`�����{����S� zB�QD#�:��zJ���/��D�A*#��ue�� �b(dg�2:ڬ����~���.�59ك�ԀS�r���'����k}�I��Z�#�Lf��}�շѢ�e�T �A 9MWu���0��%�}�@}}�Pk�y�a
]:u���R��?䵄u����O3~�Ҙm��P�9Lÿ�'ɑ��B��ﲺ�@�N�5:�v
���㱨�P� }#�+["��<��__y���0��i�<��@Z]�n���N��TWC)�	���˽�|j
�a�X�k�#N4'��<�����C�	x]D��h/�K�هC�7:ܛ�����=A��l��u� �L:���)kS�6��y�`�JU�&�P��I׷C���m�;�j�߬�YԺ�e��Y"M���}K���X_ج��|ǜ`x�c�n/������w�a��ʋ$qׄ�CmJ������ykپ�DHI�Qu��CI_!+c�p�ϽΩ�~�3dXa(��a>�J���S2X6ZU�!�k��:W6�nck%&�t�{��}}���
��#Ҹa{�DtQ��S�r_�۹�
c��A
njm���I��X@]L{
xy���`cح�T�W>��M)��}���h1T�CC;�t;���9΍Y9 h�<�tF�fB�F'<AR�|�����w���*/]��*��zMLt��P~~ւ��K�P�c h|�ۺ��Q�{8�hƇ VI&B�����X�ж깃�%��Y�H2�t][�O�4F�#˪�������9S[d 2Fݞkv�ɓ�az�͕��P�O��Sx��l,��Iʹ�*�Y�xy,wk�y�Z���l	+'M��+/��7��ۆ�������)A�iz�7�Ob5�!}��T8!�w6��[n��O��,�4Kn����I��2~�ps�u�1!�s�@��R�>�
�QK������a����͕8e-voBc�������:ȳ}�	lm	~�θhU��OFA�"�묫�4;�d9�l��i ����e痴��[�HU��1�����?v@���`�������F*�4�4�i�,�=���+����b�L�5au��Ή\nk�9ҽ>Q?r��7�)o9<hL��n��#�77�1p8]q�pȔ(E{�~����6�����_5�p��"�H�ǬeVF�nQ|��]�^>�T\?z 4�.�\�������~>���5eV.=�z�L�qXf:�ɮn��R�z�F������c���l+#���@vC�`R��?���u�v�.���:�k'��������Ͻ�m��p:;Z�V�vpj�l� R )��!��{�����`/C{ȡ�ӻ�ٚ�
~��3�/]>3�[S��������n����O�J�m��Ԝ�Gif{�����j��i"�ڟo�ȵpF���.���sp���qZ׃���O,�_��ޡpeƹ��q�,�w[�\� �;(����ޓ�_�[��0��-
����TD�'l��{Ȓ�<�a7�.�,դ=!��C�P�H�ϫ�t�r�[3>vo�	;f��N:2����X�\=��x�d��sL�&'1ҺB�X}(_3�}��-F�_����x�:�PY��\K�uî�)��7��� .%,�������l�7�(<ݹ7j����K^u�\\��)z����dҩ$D˾�W��6/9:u�,>vQ��ޅ�ܐNMA�(�R��)/�K�,�j���#<8l u��:0<��֑�P��q�[g;�A&DEE��\SV�/
7/#�ũ{�����ixnh�	@H�o@�h���~���c�B�~%��ϟ�h�󗂡�Tgy�Ux�v�� ;�6�n���c�wk�E���D�tc��e��,=�Ƭ5S֪֢�m-�)ן�ܓ=�� ~]Wp�uZǪ�|���,����l5a��p����ۉĹpklT�r��+ҴQ�G~�0	P�M�cs��we���kry�O�����1i�%��@�}U�)͍{~��P��5p�m��yt?y�)��bZ�EO/!vP���3l��:���
�6bC�msk�0��޽���hay�;�s��IV,��#-i��݀䄣�Y�㍙�8Y��i]I�|�	�j�r��o�7
�f���JyW�
������_r��<_�������+�k܂�,u��d��q��c J*?�iX_5�����1��S�C�#x�{�;B�슂�I<���XX<P�Y}��CO�B��ku�ɑ�p�9rh�����i�Gբ�*������+댥sO<���x��tL=���_� �w���xb͆T����4K����N�9)LwxS�]C\�n;�W�|l9G���d0�(�����O?������Uw�ƪmz���F���]<��x�n�ުw��,Q�7a�;�]��)_�z�&ۿ̨v��4D��Fg�4X��@M�D�6�u����|�x_~Ϝ��l+��Y����0T$������jPeH�R�r�g�)P&�[�����G������ݕG�[倽����^�kN���@�qt���85*��~.��
ʜ��F�V�De-l��.� e��X��((ME[L�kzՅ�Dj��<�K�/�����3��`ق��B�������f�Z�;���XGA���|���I .��G�<�>6}�nZ6�B��!p�A���	���AMU��lR�"���ǣ�����/����`��Ǎ.x ϰ���ly���D�6 ����'�����cRt)�ݸ�ǘ��	�jK(��lv�
Ɓ�7z��ɧX�-`}��5�怼��͑%�cC%��@���NK�%����H�d����
��u4���ǠV���:��O>�?�sI�K����6Jܰ����S�ٱ�{*�.������b���R��i��G_X�k�h�u��7��G��g�!��t:����l �!)r i�$��'0-5�w�ˡ6���ȁ��b+�l.������f7{o�g��ZyG�l�s^kLw����"?�c3��6�	 � �dV�uU���O?���e���o�bL�)E_ ѠT���N�f�5�W���5�ʓكLP��'Q'XWx9V��ܘ�X���xg�>H�/��fX~Rly��=Wy�z��A'���Ö�g�J��Ǽ��!�I���yӒ������2l�y
���{��t�C�f�լ]�����[�[@��h;ά�ZC�U
DL� Kn�L�
�Ҽ�]�N��x�W.�0���`��l����gJ�a��H�[0r�x��7$
��������f�驎�v�$�?������G̻ώ�|��O�I]�#�yp�C�E٭YP�jUֿ"�Z�"��l|X�mW5������2)�&f.{����ѣ+��~������>�m�n�1D�
!�Dao95�=��ؘ�h|�2���hD1�Q��[�!�u&�M�DӖhw�`�Ǣ��Y7�����(>�:N�;�w�F�6�j�]C5�ǡf�v��f�Ǧ�t+1� sG��\ĸtu�6jL�(�͡
�����>���%�\�*ܵ'�1h������Rb5�#����V�v�p���Ĕ��e��R�&6���������7��W�1D�����N���Gc��	^�!C��֜����V���O��,�e���>�#-w~Ĝ�FVO�g�oܯO5(��q&�D�+�t�f�Y����S�/�����?i{j���>��yP�q5�&J�w���p��7qJ2�K�I������Ȫ��<rןd��C	�&Hg��BA|5i��+ɬ�Ҕ��� ���/�[Y����%�	�3>^l�#�dKR�x���q�	X�_�oc��Vy�2���"8/�<�������T�ݟ����L���]ɮ����E�p�e��2��l����a΂� �X0膥��X�c��/ۚk���L�h��LR�WIʧ� 
��_�=gA �7�2�� 2{���Gc���x����J6��F%��c�Bm��b���;I´m��Jt�E<PiȰ e��Wc�y�Kc��%�M����[F��h;�@f��l�F_>��H�-��V�R�mO�����0yD�{}��H�x�0}#Ǳ�^Ї?�8�Bũ�3�Ѷ����.ء̣A�?���L�9^�g��Z{�P�i�^�I(��՝�هm���3�vk�T�O���"��P���������_��"e|=��^��ڥN�H5�6QR�`4ZI���F��5B��~��W�R�MH�W�gG^8ͫc5Վ�5[d=�TW<𵽊�ۦ�E4��2�r��ny끐Zԣ�O5���(��·�
���{�[���-�)m�Y���˹Az��;	�ryWe�}���@U�/���z
�)�(�ʰ��F�s��"_���܃�$�CjEP#�����٥)�A{\�x��� �Pp�:F=������$Ds����)^ë�M��ѳ�d!j��F�6�Ki��z{E��GY�w�v� =|�Li��L�e�Lm4Sվ+����/�?(�� kGv���Dɀ?=��4@�������=?
�ir_�/H��E���!�^�j(2T�˓~��;���B��1R�	ԦW�� �ݯ�j	���_��?W��9{&�V�kѣ�T�͖�i����+|��1tٲeU�ϋ�M��q$�?�♻�~=9��O��?>6P3
8ٝ5_����	&�^|��שS[*Q��Ը@諩����9I��ͻ�w��cI��̵5�ٙ���U.=��q�?u�8�hE����3r�Z��Z�(���������l�p*2o�Plt��7��t#�f�ޒ��b�l4�aŻ5�h���`���e��s7$�_���\�nes��Yءp�m�e֛�����ច�b<���G[��,^��P�"�L߳
�)_�P��j�W����P��F�2.���F�z�.���l-Rkq�eXm��ͫ�2+(�%��P,��+$�=�=��#l?/�!���ƝZ%������A������D�[܂���I��n��x9gn��Q@�=8BA���1]�&�����
EAѻ<��}�z�[E���;�7
�w�s�ס6R��d���&��P�LʰNm�>�v��e΀ĺ���1��@7ox ����+�n�RZ�ȡU�6]���&�v>}�7�����{���S)Q�Q���o^� 
�����1�v˵� (Å�x]۳����
��|a]mfE�h\��;e��,�̅w���|���ד��V�U �	��~^1�k�`�����[��v��l�����,��p�\ ���A�wq��99�l��.�t� ���ky��ο���Ro;�B¥��i4Sd6����U/�)�7��PK�r��$�W�QO�cʜ�Hd��W���9��d�yxEܽ>J�i�O��ylfl0�~���p��ѽ�׾�|-��s�j�\>\9	�F�ӗW�� W�����H��YU��f�t�|e ���.	�Xi��Ԋ�� ������$C�5I�Ć�=��eJ���ƥ�Ξ�n������,���������kAlL�q��� l�5�R�t�ɿS6��.4�
�t���f�ޞO�J-��]�3	^�Q̹�'��̵<p ��(+$��B��_^�m4qe��-K��� �l_����nC�/[�¢:��H�J�w9���߃��s7n�|2R���	}k���/_�7["H省/�TBƹX�Q���ۉ$�7��v��E�Q	j�.�u��0�
�P���ū���(1�ķ���-�vK��x@i1�]?ή��$E=%=�1�]�_ ��G�T��z��4ig΍��<׽���_��@�r�����=x�AԶ�\�U�ZC�`��+`�ְ �<Nu��vZ����*�H�l�)�o<9?�?d/�c�ĸ�Go�ɧxR�ai<��8��� �6G����:���: �BМ��vPe�f�Q�+�Qh�`q��B9�O-�{���ݹ�L����-=K'�f���p!�ݶ4�4�=� �N}G/����ynT9��	����p�y�L8���"9�+����&P�⍱���d_�Z��X�4
:�^�n��6�|F^�"�0�ceW�_�?w��J��-����������ӝ�`��f>lz�b�v��w����V���$O��G�n�H��}��p1�d
��o��!����ɵ����)��4�._����A$�邢� ����j�
uj���{��Aӭ�X�2]����؂�Z<�gn۲e�k��f������C���� �
�7��>�h2��r�P~r��=Q���w*hPnW��á0��%�޻bWʹ9�AH�zx���7�6�9�ۇ� į�e�$�<L^Dg��5��g� ;|�n݇��$N�{sWF�x�Ѳs���'T>��ʇ��r��DS^�Ic�W*�T!,*�7k&�Mpφ���N�ΣrO�f���CO+��ǰZ����u�,�~�l���e���I<uҧ+��<{�#��#�t$I��2 ���w�~�����1����v�Ҝ�ƪ��.��1\e[L�`{�j�k�B���M�2L��>�"�卻����v�D9	����<�� hH{^eo�|);u
�~	��s���x
����W��bϘ�`�N �# �i�\L|�`�'�vXZS�7��^T�W�,?���)\jU)#�4y�R��/�I�
s��f��p`�Ӥ��U�=0��U�`[�i�|����v+Yn�J+���P6�!<��&���0ξ�ﮊv�C�"Q�^�!�sFϢ���	��vP�C�gf'qgť/��d]h�u2�K��
�Zj�P�� ��V�X 4Y�z�b<C���ɝ��j�˔����|��z�y9�r�Tu6�x6���(��&<�eo�w>�謌���v�1j��i���K�n��܄�w�FD�Ʃ;�&�nő8�WD�L��7��qڎ�ۅ���S)X���p��'$�p��e�"ƋW�_2���ov�V��}��������_��f���^E� TM+%��O�u ���r���&U�/0WL�n�(�F���0e��j��?�Z�(���Zox���A.�c�|=�Y�%���x.�e.p�(��я2�l�kǧ16O4A���0D��w�B�''j�k>�[��)䳂��@�b@��t'� (��x��!ҡ��+X�L�3�d��	�J^IV&k-Ơ����V�X�Г�
�4��g�W����x O�/��`)7�{��Z�4��������ËT<q_A��}�E7��.��-���GIJ$nV��I�Z���!�wD �j�~Ħ՝��������sA`	���l �={��J)���zRc�fX>Mx�(�l�mj�x<GSqj��{ ���Y��N�$x�����`c�:.�WQ�(-�V����e	�I�h�׆����O��5�P��6�n�WX��ή�$0��oZ��y�O�ۄ$j��{��-F�r�}g@9<�Enm)/�'�3�[�ќ��B��W��z��NS�.|�����9Y�/B�&Q��^B!��ʊ��D��$R=��B�Ԡ����,�-�_�燡�-.��\���18����4 >H^0��yTj<C�R-��Е]�!��pG���j���5�8hD����
���_4��?�vH����M o��*��s�
<zB�
Y6��J)�D$	�bN��⳧a��F@eW��6Ø��/{��UE���� Vf5:� S��M�5��4���n��I څGp%���I�x.��9e��?��@u3����jF�'�Q
�؜��U�v�+Ԭa8�Ȓ���\By�� �q�\�{���+j�p�Z���Y��w����ţ�%�4̻�+D�����*	w&6o����qx��W���Q��X��� �R*^kO�x��X��އ,��!	 �8�i�}�¶��g�����c���Z�J�'��]��plߺ�1
*�JoMB��Xͨ�{f���u�(2��֜��Y��TR�z �:��A+�IK��/�Z�<M��{�Ѡ �f?�Z��s���*�o��\�=h�dܧhb�z�j����P��ƫ����`5F��y��b��b������(|�SeȤu�1������-&V�_1�體?$�R��Yv�:��^�۽�+ӛT'Ͼ�&���\��S�~�Y�����]��ԴpW�!O���]��L͖��7� �,K���9��남��Z��'Ǘ��&Ф�,�a/ag��@}�!��|.
Yt��N ���j��ę�=u���a[q5ǥ9��l`R��Li�b�PL�����g����`��崮�{jPG=4����<����g�g���&o�n�:��2A|��o��U����=z���o�~�N���y���d85�FЬ�VS�FaG��D:p�)�;)�l�Wb#ɦ��6V��#�v��E�*P�eeņC�e�!�?B�����q�My����E*�K�t��S{���1/�#�!��ۙD|Ly����'�.�|��Ѓ־���"����ރM��GL��l�
2bY�u�w���{���
ta+>%�#khk��bDԙ��G����j��g R V�0��7�e�ΓQإ�����'���p��cI�7�H������?'��C�2c�"��qwC#���]eR� ��g?g�1����-���U�*Z��q�L��~*,5V�_(�R*�K|�I՝�s����:u�s�㹨A��y�p}����+��-���v�����Na�Pߛ�"«w��՞Q�X�o�]�Hӑ��#
��Dw\�:9��*�3���J��'���iH�7]"l��#�x</>ݹ7�	r�Q��ߩ��N�a���K�<�ת�9�I�$%�G���DEE[(M�4��E���'9>��5G�W�m�)P��x���&�|�������J�{�,?2�s!�a7����7��n����29M����B���ye�mQ?�9�.����i��cU(�\c�����r�� B��@4�K{�e�/����[a����W���f	�ܠ~�g򪅘����Y-а�=���X�H���g۩�0Y /.�*'ܖO`.�����������Q�V���������a�ۛMʤv"�qrb��^�5�_��q��i�@������BE�E?
�ד=��|Ye��p��M�S���^��9�;��݈��7�l�@,��ܿ�^͟Q��܂	��y��D_�3<-�hp�<g<���Y����]hk���%boYwW{�a%��,���h{n^����s쐦�L1�����ĸ�n���o���l���K;� �i�`��Ug��O�~���r,���Ͻ�=N��\�w�GÍ�݇�s��S���Z� ����p��Y�ݖSN�'U���p��^9�ݣ~=�s��g���h�����By�1��b6T{��kb���;6��WF����LCϞ��IYi�j���{��'1�\�ٿ��[��m� ��Wr%U���0���a����e���J~A�����1	�R��us*¾��
�;Gā|�~5���Wĺ�'��l�V��19`c�~k�O�\�h>:��6<�	�ӰQ����"2&ұ_ӳ(fp�	�;\�؀�|x�e_�����N7�{Z��K��^ �u8d��M�1�δ�����&iX�M��3�%eM��������~U�P�	��Q��!��%�3o��΃� $�,� υ�d�B�l"��839ҕF��
V9+���?#�'9ߒ�I�����E�q¯���b�(����oH%4�1���,��k���|R��=�=�3^d�-�l޽;}� K��x��+��*o8�f�(Ys۶�]X���"��=�N{ty��u��oM]��I��
����V��{j��jf�+��٦_�Y?x�Sx5�sׅ�X�;x��)V��{��j�yDZ���&u���,j��Ǥc�����I�#��Ң17��D:t-�Pk�'�,�b	k��o����=�z���}�t�����9^\�Z'��A~rp`��T�� w9�����@�5�7��Y�`�O�.����|�(C����Vp΍���\�B:c���Vd���x��-�;8�uY��@M2�9ó�uh�J�b��B���Nou�#�R�kk�'/��؏W���M������L޻�*��&�Km�|Ķ)][��Dy�_|��.�H��x��=9�j���(;��=��:՝jo�`v������pě|<V�f4��mY��jy��u1� �ɥ�,�G�f�)�T@.��1�g:��(ɽ���։ ^��-5�`�xfG�D�W����Pj�K�13?����4G��;�����i��8�MfӷL��H��c,ob����#y�#xW�E���j���;���6�1�/��#�	z��0�EV����XM5?zÐ�m$:k~�i��8�a����s�G���^Б'x�LO�ms0����#'�t��,�v֋���cԏѺ/���&��WO���4gσ�7:������������Ba����(��@��C(��׮�r�8�M l5r����D*��'U��._��uιo�f���ƶC�v�cц ��@�d�H��>ȿ�oAD�8:�ra��~/a�On�^�osC���H�N������T9�>w��[�-r7���@S̉dъZ�3�vj�Ӻ�m��D�=��=����ZxY�$�RV����R��dXnGG^>v�5���ο�x�ќ�F��2a���J�0�پ��U
��j�J��R���>�� O|�e�;^�b��ɱ/�ߵ��KX��E`ru_� ���M�<��ƛ����)aeg��Ը�	���$P)�a= U��Ҏ�o���i��M�v�|��{�[YQH���t��n/�i���<��S��S���n�=� @�p<%T'� 6���ɡ��TPϟ�P[�l��0���۴sX+��ZB�5����-���{�i#u����t���Xa�����dL�֐���R:^@�n\�cq�P��s+��w#l�1=�P �>Ť���E�9�a�3l-�t+z�!m�)��И�OR����p�-�[N�{��-���i�Hn��ֆ��p��Ȟ�j�S����t��-n9�����,(�??��f��]M���[�89�Rt��h�4yc����ILY�5!
*׳u&�z˚��x��g�n�X�"�or�)���u����(�$�QQ�e��!±ȹ���ڔs�_HaQ�����M���;V�ʒ�O��+������M�z���5|!e"��;9*��s�$��-� �Dؑ��zɜ��ʦ\�(��Uj�P�����V����� (��Z�� �i��F�G5ow�g�B(�3X�e����5��\��RE(a �8�[|�7��`v�x>��~�GH���x�����B��B�dQZ>V��9�����w�S��1R��4L�|���p�(D� ���ռ����B/-���<����%�1|QF�����F�\��/��8�i�^���Y�,��>Խ"ov��C�M�#7����"���U^�<�(�Ww�6}G��� 
,N=����5#�Tt�o��4�
�L��2�Wh_X���T���en�r)���
�}yY�o����[ϻ��A�Й�d
�f;���b� �|�np�>k�p"(����w��ˉ̓R�M�΀b�p�\D^��@��H�9��ٶų�ntb����ks ��2�� �$�u�&��u7����_H7k���%�>8�������_��x"+n8��gV>�R��{��K|v��&>.�����M�M�o��ﱃ��m���9 ��PQAW��K|�^�/(z���9���"�%�����?uz+��3�%����]��/i��ѥ�ү��?]���9����/�=nP��/�3]�S����gR�k7[ .��;����X���;�E^�]f�}��ߖ=���Q�rB;_�%� Գ.�D�����O��JR^2=��KȘ��u��`g��jg����%�_�?�Ui���{y&G�͗�Ʉ����b=�9�����::�UR^1��m>qJza�T���7�b��.�-䜺����CB+�p����v;$�4;c�%}D-�9���~�Q�@���� 4$��r��"6���&�{B�Rdw{٭�~$����6�t]7�c��.D %���d��JUq�e��� :*7�&crŕ����{�G��d4�����0���C�a�-^��"g8����G����&�Ϳ&�K�n��E%0ި�с/d?�ۃ�GPny�Z��
~:�N|�W{���wC�yQ�3�1��P�U��E/�ޓ��s@���	k�}�z�F&=�}C�_���w"k���K5��\/�~�P�� �ſ��ȯ����@/�b��+�K�<������23�13�13�13�13�13�13�13�13�13�13�13�13�1�a#����,���@���@�󘁍ؘ��ؘ��ؘ��ؘ��ؘ��ؘ��ؘ��ؘ��ؘ��ؘ��ؘ��ؘ�����>l�Z����,���@���@��Bf`c6f`c6f`c6f`c6f`c6f`c6>
[�d����/UEp�\�*�E
�"l3���$�pV�'�w�O����:I�s"�.� �M���b{~�+~6*�U��8:�'���ȣ)#������y����)��#��d7OR`�L/�򘔧�X�_�~�g-�`R�M�$x�N�F��8��j��})w��Pw|'����듯dK����G)~~�c��i.7R�]Զ������ra���-Ni�lU��;|�(b�����1D-]��܎G;v]X1��sW�>7�g�:�x���I �z	S���e:�ԯ�Н<Ӭél��G�t�a�<�;�	��2�tоu�Z����??��.&��;�U,^�������9Ca����X�c�5��P�]��=�%t����QY!��[ ��b�c�P�N3:�lA����n;�زS��/^���Ҿ:F�4��<��e��տݏӑ��!�7#��3��$]�DY�� ��G�ˣc��O|�&'�ð'z�J�LZ�HWe�&�xqSs�m��>u��⑼M���s��
%<�ḽ���3$Ze�y�wgΜ	�����D��ާ�ç:����4N���1�?Y���K�{t_��9r�'z��!RJ�Sd5���A?�Fs6nW{m��6�\2�>FJ0_��&���#������,�-"��/�1$}ly�!�4��]X�`>�/��R ��ܔ��o�J����:��p(��*VX����?�)Cvn���2�h��>�<N��}���4h>��kfq���Z��bp��=9N,ߵu�!N�b^�H<�^���#�p�����䴪�"YRw��͈A9�SJ���
~�����9��_��f�3�>����7N�p���G��w0Ŝ[=w���{8��.�h�!���s+��`�p=&F*�J=i%p��7ꤋ��e^��?n$&��,�OWs~��xC�����n��+�~|d�|xb��RGvǓ���	a:�jo�눻�$�{W��c�=�U��};�e���3�ҏR��z��+>-v>�j� �[� �x���Y��@]�G�G��S�Oq{�c������I�X���܍\���r�������I�\|�=y�v'����6��D���ʯC[�	���_�_� ��v||��Ꮂ;'�S���|��`�֜��t����u�O�6�Ǣ��~p�57&w��ǆ᧔�����j�[��~x��%ߴ7f�8��>��To�V�/�cOo��|*Fs�%�:����l���1��akC�d���Ҷ��8�eBA�&�� y���:��$�XA��v��$��g�u���|i4�Dɨ�����ܩ1s���X����m++�S� �I��;�ze'�/;6GT�Y~��� K���h��Q�oe�����;���jи��t-�1���r��e"[��H��egX���)���f���5�oY�����'�)��zM�J���%��{����N�v&�G�E�)j�~(��V�g�W����_[��?�����}��.6[��4/�`���c���Ӓ���$��Q.�:�����n�	F{r�c�S��~ ��/}�Zu�uC����...	쯿�Z�t�\y�؁>�-̟�9(�8�9�n;k��H�4N�1�����ߺu�im�r�
��&I����K�_Q1���c�ܬ벷Y��c筒�l���/{����Ԍޚ�KI���5'ӑF7��3��KS��
~�z����W�ŠM�_۲r�����?9�S%�̣��ą��>���� HmA}��D{���>�y��_�
�$��G�Z�ƨ[eT��n���$� jd�\/,{�4�u���8#H���Xי}�����:�jYY��d�ԿO�>��aUd^�.���&�$QZG?�2xY�s��e��7��}^Ք�TZ�d������,q6	������[��<q �G*#���>3008&����w��xʋ�ܻ*�l^=��}5xNǘ!Ͽ���>�K�&����V
w�a� ����`��f�_^g����_s���᱾�k��W1M�NN�ϝ;W��H���K���,S�g$폝w�P'^UU��^�ǫѓO�;�z(!���޺�w�����mL����"���$e�!J��폔�E�wO�8�ix^���4�_��/lʦ3��o1Li�sL�W������D�|s�pc��~f�,@���
o�H�q4�2��xrҩ�9:�=)TDDdÂ�'4�%��Ȝ9��)��z.�|$Ӣ��R�g�֙W��<y}��ڈ�w���~��zy{{����X(p�4ʕ*6���dd���`��]*�����O�Ք��;�7I���R?U��+�W4�1�b�^�ݟ� �ה���܇z��1������iG�I����X����q�(����jT?���)��ۯS�����8�f�����9�J�u�[��D=�\��9������=���A�`s�:D��ē^-D�Uc"���x�=LFm���X�܏��V�Л�wK�g����$��˅Ol�"�I�lۺ5����^̚=[t[�'�Y���q�U�mw+z���������m�$�U
V�:��Χ55�"6��gfM��|^���<��l��ĩ��̓g�̓mc5<O��V���L�c��BX����jP+fۺ�1ssӒqA��?�y��L����o���,��	�Ѿ�������H��BP[�u;�P�}��\WA`��J���(e�VYNɑ�x�`�O�^��3�wY�Z���њM�5��ܧ�*˶r�bwUt�z�ߺЫ�M^R�z��P�f�=8�r��:���HF(1_&��T�|�ɑ���)��ғf��P��EmnnFN,�o�[�{��o���84�*����Ð�{Q*���1�C[��?j����?R�u�������v~���W;�*�uv�8�*oWe~�?�t�t�jd�Tb��b���,^�]�Iꫴ $)�ȱ��v>�o��a�a���cgݝ��{�����J"!r���R���՟�g�R>=:��aR+��/C��V\]�^D'ίO.�~�k2_�z�N6"-u\Zr�a�y�g��yL�	��a	3��a�b��՚�񗏯ͫ��f�C	�-w�e�)H��2���KRL����>��z������Ǔ��#���ց`��A[dR��Z�"?�?�ӹ�r��5���M����:ztۙ(�s���Y�foSQ	���
 Uyo�c~�ue{S���P�o^U����#s{���l߾��D	`�C�;���>�l_PP`��������Ѕoo�P=�Aє�w`���Xt�-�[H?�Qe^ّ�'�jc^/m���Гg[�0軞4�d��cj�=4|��o�����p�������9����uQW[�eg+?H{bد\��֔���؍J�@ze@��Rv�e�<tU���� �z|��r�P/)�����h��Ա	7�h��h�f��j;��^���'��=����Ts��%!er�K���^�7|���ᇽ�*��u8���2Vԥ��Z��%
�tt)(hA���H��0G[\L,PZ����f�?#���ۃ��M�������h����;謺ZLF@�����#w���3���R�'������o��-WG�ό�{�p��݈�]{V���'b�		�$?i��m�QP����P�U*�,�W���5�|�c~�>~���0��"��r������6�e�.j�RZK�U)JOW]�`o4���8��k��=ձ� ����-�汙=�_�A��rSc�ƽE^����yʏt�6��'��C� x��z�,���� ���Y?�y��2�|6\�z��׎��'��쓇sO�<'��'ƛ�t��ܒ��iG�<xY ^k}��κ��j���hl��fQ7��1�R�cccW�U�ikN^�/ q��<0܉���=�FF�y��,����W�o�cӘe���-�E�HgEE�x<^��2�C^�,G�tO���K��N'��b�~D ܬغ�w'�8��wd�6��u��x-Us�Q���� ��b�2}���<.�����w�qNT��8��HJ5�#���}D#i�^��P9DH�:R�VI�uRH�j�Ni�SM�4��z�Xo�y��~���u��i�z]���xޟ�kyё�eހ����%�5sLOM��r{����k7��ھ��r��4����YI  �t�[d�V%��,g�=[� ���K��<�Eվ��iH��フ1C%4IQ|��ϼ�7ޛ*ҵc�|O�'!�M1�;W�=�U�*�F��'Vt��B�����d;�~��^���W��wb��}N���CC*�j�V�������ٙ�~���?�ژ�n?�1��#3B�q�z)�(Hݸq#�o/	�EW5��%"������-�=���<�OM? �⃛\6���}�[M9\�޿�Ĝ5��YN�h�"�3�2$Fi��꟦���&��֐�����ck��'O.�o��1�4�B4J5���/513����?��+�IG�{�Ljlj�@���*.�\Sa�2ś�mD�ezC�{=6��ȡQ����G�l�+(��3���I�dM��A#]]]�4U�j��Ё�}-�cG���z���D���V�$�ޱ�U�b���f�38V���M�=Ӈ�{i�"��}�ao��<O*��@8Z�8+i�*��h�5߷ ���Q��*�j��@c'��b4H�!_w{��o���X�!yШ�8������m�]f�E�jH:M�M�����v^� �ɾ>���@7T���g���q<>���Uj
�s])�p���|�\O�ڲ�宙��a�q���VVVs�ܧ����"����.�[F(o��p ��YIw.��_��%�����7{<>��\b4l�	h��8�;̮&n��b��
�f�I�4s���Uyv�ٽ�U�Ĳ�f�}����;�ic>��p�V)�l+�-�J�#��י�6�j�2���@S(GqI�CS����Sk~"���y݊ʦ�h^�����/�	���l2�b82t����Ɩ��9x�9Ղn��ͥ��#��,&�y����u�]�ۃ�(1Ӟ�m[�c,T��8d���]� �lG2�(�a���j"�@ӣ��GT���KCq�""�U��^��\*��㞱�RV��m'�멶G���B�5#�ٷ�{�N�e�aV�iU�^-l�<�����W*��L�;�olSP~����>]�!s�b��݁�r�ͣe�	�(֥����BzQ`v�uy�!@������٣�[ ��:3�:�ks�����ϟ�����s�qg���Ӄ��yZM̸��G�N����2LX�G����B�9{��ؔ�?CĀ4��r3.�/Ȁ͠��ѭs\�>H*D!~��hϳ� J�@8�~��׼E\s�z0tG�s��n/��mE��s.�[!��q��Ո{�NA�z�=�oq��3czko�!ryl�r��R����l��ȡ]��P����_��Q�y���f�VA)<��G2Ѣ�Q0�^������?DRS{T���ň���`����J��j_���W����1R�Ζ�#���#$�����9BF������ҧ�Ӻ=x�����<Ikݺ}���N�L{L8ޱu��ߚ�|���g�50Nͱ�t��^&+�;��ep�j�X��h'��Ʋ	F�kż��1ar�h��j�^6��xE)5�� ����\�(�����_=O�S�6�-6>3~�S�f����� �$��ުC%ׁ�oصkW�'jRbu���}@�����'���v�U�
��Հ8F�iXJ���F 7ɞ?D5�w�45.���o�r�'���[P�w���� �,#�)Y竗�䴼�d�[g3;md�f����E7����׬d{Zc�]��y3����.0�Qdrl ����@_m~������z����V����KZ<�\������l��B����{�Em詮ܖ�#�� 1>D:�oq�ջ9X a�Q�@ir��Č��g5VWW�J��ͽ�G�Ҿ2��z	 .�
�-�UGw�	Z�x|�I&�F���D�1�M�����o�z'�;GJz��e�oR͚E��_L��	/T�ԝ17��"�w>n����W�J�fP����� \����`�ᘑ[D����I������vP����t=��Tvl�����|�n����}�*Lԡ����E��[g�!�ny�l�sXo�u_c�I��;|h[+��W��)���0e���I.g������2�:sVy�*v���eD�K��6IKK�|�d�T`�a���qN��tU�QR�h�$���O�칺��|�ד��X��M|�c��:�͘!��I㕐�a��`;����x�D�v���I�/����ݑ�9Z��@�i�4���DJoK?h��58�;��<���+G�Z����Gb��.<Xtw������O;]3�i����W�2���"_!U��� Ӑ�[���-uus���*n�F?[�w��%���m��L{��E����Z��q��3T"L��SdvFi��Ϝi|�p�f�o��U����A��(�����s��4�i���`0о��\����nRkk�����uK>�C���;7%e�ic?�_����N�Ɛ���U��@�V�d�|N*�-�j%ms=�"ؽvS�ΰ�+r_�1��F��|f	-tn�(��!F�-M��]
��G~��#������W��Z�wG"�wi�˙�n6hc��#O��[�N�"��vG���Z'���L��ko>��w����ΗsK�"�?*H�r���1`��=�	e�T���^<<��Qf�o�<G�֟ˍ�e�@ef/����>(�n�eR�C��I��)H@
U�RO��9H���y:��ĽM��\�q�%������6����R��b�~��� k@��9��ʺÕ��A���+�f�:T��VNK_��f�����t�D�\���T�V�=�Z��i���g7��
��|7�N(�d	�)��T�"W�Ɖ���V z��͛'����}gS�]W����޽�G�}�L�:@����>������[�c��@ �i51+�y��= �a=�t�át��c U]5) ׸��%Q���Ë�4J�i�6����އK����4�V�|<�:�Yv`�13�����$�G��捷��(�k��RӶ��G�ήe�̬���D�;3�O���E�@��y#j�ɫ�ԡ���Ǖ������MLL.�̜9���?�A�d�H����7��u�p �ζ�K�cY8^J�����^�Q�mV�PD=�Ba�Ξ1h���x��#O"={f�F�כ���)p�Q���{v��Я���
ًQ(����8}���㮮�Ж$�+jN��D�;H!�FY�s^�S=�_ "ȹ���MM�>��;Q����L�sl���Q�[4_���C0s#Տ��D:���4�!�Fؘ�J���2��������,l�����ٹm>���2 ħ՗����N�bx#�8�:���˳�෇L��$W:�/����]a�R�O6��F]`�aA�,<#1�f�2˽�>Ѫ�O:�X��H���UY�	[�:3��Q@Jz�i����cd�f\�����*w݃d.��nX��]��Ǎ(M�ep0II
�X�mCIB'�)]��pGi H�t�7�H���K��F��aUd{/t)6��8��"1Ʋ�VF�j���ի�[��3:>�a��o�_
�� �3�x�U�k���
�Z��Di2�{�9��؀<2כf;������ل����Pw'�(���;ڟ���?)�4{Euց��O!]��Ikkt��*��bB^^^/)�h��C��tŵ�� ۑ���z��*AN�s
d'ff�BgJ���ϱ�7
��R��{��44�X�(D}�l��Dd��O�u�	_�`bn:���PD�+I�c�������������ʐ���� G��8���E|�����������9�#nG����/#����ָ?�i�������{=��2v��
���c��v�nL�y�鵩���m
2����4��|���2�q0�%�6�;�!H�c�abu�xoC�X��v�H�V5����x̘Y�D͙��s�E�!�wi�"X���\���HIgYp0��m^��s�܎�j_5�.Gf���cXn�מ*8k��4?29�]�iv���^��қ��Zt0d�-�tK��U��#���V���;F���(��Ψ*X�@5y�*�Ֆ��*��tzj�'��P?�_ao&$��uUy�������w���Kx*#"��y�NJO�G4��
Gm��4˜_�펼�&�ڵ�<֭R��g�~�	|M��։��ڀ-g������������e<�$@%�[!�N�=n{0��][4�޹���V����F �r�J.�ِ�8�H*���P�Q~�Dk�2I#~��X�ê �t��3�W���q�@S(�Bs� v�v�fee-�w�zvo���]]���p��Y��l�Sk$ZI3y3 {E����B�`�-]�lw�HW�t*�5z�����y���(�`
3C����ռd#��(��e�>*_uk>�mW����к-ӟrc�Tt�@��OI�@%ȍv{����>����v)x�>U���Zs7;�ԥ����	V�QTblAsLM��Ջ��m	����l��d������)9�ǶPw���=%�� ���{CL�����͐��Tn��y���l�ӷl���_`eeeP-�uj>eN���WG�3�q9|���VR�-�~����b�K�S,J�U�Q�)�ʫ������/��Y��H3���s���-eE�\lI���T�C1R
�wl�ԇ���m�aG�8	?�qu�3���N���'��M9;�+$r=RSl���\��F��
����`^rN���F 5v��ߖ�?<O��`�ċiz�O��騏�����%�4�D�Ĳ%�Oor",�J��W��X�dTz~�^a0�6Q[�;J�s�A��p�fm\6Y�P6��W���˗���*;�(D�H�B{M���Ĝ*��1�[D��0 �G(D^�9Ֆ�@����������ώ�������Qk�B�3P��ه�{�`:Ĕh����]�dGq�1������=��*BL�}i�z:2'���(����a��W.p^r:��b6��,p�쾺�n�JP�=��0j��3���}K�Hi��OV���9 \̟���j�L������D�\n^��*t���d�q~�= ���ħ55{}�6&�*�Kh5�`�`�J����.;p�`����jZ�,.oh��L�Az�Ò�G-�@K��Ԟ1o޼�\�[�ք�a�r%������z��π6��K2N�4eP��H%��^|H�G�q�Lo��&b�bB~���H��gy�5\*��B�F\Mj�W�]���J�����Ԍ�kPSU]J>阼g�%J�{m�|�T[6�=�k͇�鈆�0Ω��cdMb!����gi�n�YOl^A�G9m�������7���=U���>:7_�~tf�Y)%�r��@�̗=�d�I�Э�����q��/F�4f*��ą�������������(�ԩ���6*B%�=0��C�7�2.�A���fzӺ;����F�]��*�trr�M~ Z,�R��4J@����y=��z8N(��>Wڋ���v��ʪA�7�8������I�ŁBe��t&M5�a�lj���l����qp؅�r�q�K�3��?щ\���q��,�{����g����`��H�<T�ǆ~7�$�1� �t��S�����*#��-�i�a��d]��r��L�ߩ�ZHު���= Б�{.];V��؄�����'kTRbbb�(���3�^IfT�o����4�����v���QÇ���`���l�>�5��i~�hӏ��镎�Q
���h��~w����:�WFD���s��l[gjj�<)�ڝ�$;���H�-W5=M���g ��q<�=O����q�s���H{��r"k��̺{���s��LF�b���pc�2�H*=;[�Ab?᷽����}�ob(�({T��������a��l�7$^/8TvI���ӳb ќ��*�(VC� ������5O**b�u�Rhi��eb���0��� ғ���R=�!�l�--D���K���\�A���l��r��=U�-Kz~��l`|U���!`�~�&s7�ۋ��6�����&Mj�af_�˗�]�A�'G�����쏟�,��ęRۖ|�7�q� _b�7vNW���Ǥ�❒�SV���a�@'QW\e?O�i�.�x�ޘi����w��\-��N�O�����L	S>��22���cFZ8��e6ƪ��ʗ~�%���P6G�x�J-�{%��l�ȃ��ߋ�pn�x��P���Q��9]�LR-�Э>n��


Fs֩�K'�ލ�����@ȃv�\ɴ'm�P
%jW�� ��x!�g ��cs�+0kl5Y�jՁ�,�텮������#�>�*������ש�n!����9H�RF��E5ڧ��x�bYl�D��Fi1o�ڦ�0�2�
�౑�Q=e��轡0e�Y[u�f_}�����b��; O���;Oڢ4=��:v�н���w5ge���mۼ����$#���X@(zج��������S�W+cX����I,8��ǎ�����)N:�)Rc�����S�H���3@2��,�b{ϓ�G��[��w���)�2��V,�!o,om��óR����$�@L�s��e����Gon��K2	��e���0tv��Y��l0�è�_���U4GjK� ��hf(fg��U�3fi55��۸�J0d�[Bۓ����"�
�\�2@RQfǍID��;��+W���ߺuk����d�ɣ�XYm���$?����lrv�*Q���]�0f566�d/ۯi�D��H)E�Y��-�UGiM(���|��ˡ+/�59vao䏂;v�+���VO&xAc��A�d+r�?�Bc�wVV�?D� ��Gr�o&���J��i�í�����G�3h��%΃�������P���b��xY%WJuJ��B�H�R�i:�ua�?�ѦW8\��[���@ n�[�����-�(ϟ���[1��VF{gQ�����߼H����"J,�b�z�^Y���A���2�Ȗf^�D"�gĎ}Dm_��O{ɺ�����fE�Z:I_	�M�K���I�>eN҇s%�S̻
��c����!v9�$?}:��|�c�c_�E�5����J���q6��Q�[CS�>+��G���ޚ-@�޸f����5�k�fy7c��) :nh^�T�c��k��Ϛ�^�/�����	III/���W���*�խ����pb7����&1Sr��n��KWy�<��eH��et
��6k;�g�Yg|��A9f?tZ45����8����w<���'!��ȵXRpȭ����{��G�Xr���pKi:@�3���|���knp{�gW��ͣ@yR����]�������S����ڛf�*��f1`@�/_�E������(D䬏��E�������_�����)6>K���a3�AwBA��7���ݡ�DC�zq`�s�%�e\�/��6yɳo��-�fvC��y;���}r<�拾��U
b��U.GҬ����[��WA��=�$"ݣj���O~E�!v��e;�����P�ůZ�����f��Qkk%���]>u�0�ћ�����_۬6���x��Ms�XjF��]�g�{q�&Hd�Y�D<q�ǅ�x`�(TU�5h^ے�Y�g?v�Vew̢n�� ݸx�!�0��rs��pKK��)�L��'�AAw�@�ID���E�e���I�D��u��Zhᆏv��8�V\ ��'$��p���?;Xmo����kZ�����
ۗ����C�o��T�9.J\\|_~PZ!+����=rHR����ߐQ6�:�媥�|���tW�Ť��%23ttt�|��HgYٮu;#�
�9&��wGz��1�/��B˔h�sO\�+��8�|1q��tKC���Z�P���J;̺�I�9�l��~���u�(�uwYr�M��{'~/�����G�2�FU���<j1���C2$�(�cM\�\�ʯ|-�Ėt��N�|o�KvHY��3=����2$��5��x�������.�(祴��$���3w.2������ݹ<:6�tb]�Ʈ�M���5��M�O��:ZqeU���ȫ���T�툟eV�Ԋŭ��Wp8�r���Oo����q y���[�|��5���Iw�7�u�f��}�r
U�@�	8Z��Jٱ�pg�2B��&�����Z�#�`��J)sh��9Ż�6�'��8��z�á#)��]�Fr��L�Q�#hF��6jL��	��hg7���.6���&qފA�;�۟���根tR̼)�@�𕾗4E1����7���ff�'4;-#C��</>�?�}�~g�e��HOl�Ʈdz{Q�v7�ȴo�ꪡ�qў������`2��f�:/���x߆���ݬ���Ӑn�gq��V����į�\���`}��I��m�4��Mjvl,�#�y����E�C�Љ����?��]m�a��[>�����(�$�����;�nF�n�sv�ޓ����#j�f`8����è�ؑ�B�����K�+�Ewcd0RV�[Q���td�A�6_���qB��1B��d�b�a{�����e��D�c�,����B�rY��b�ĸ��r��!����ZȦ�e�a�h�?�q̐��ԡ�����eu�җ���ŋ|�\!�SK�2>�*�Kt1�*����5\�ҊP%	XG6�G%j��	��=a�{�<A��Vj��4BP3��o�q웲�{����x7{S���VE�!s
�[JV!
���9�e=@fV��	X�uk\*�1�M�����j�7�Z�A�g� rׯu�
U����ǴJ����p�A����������4
)F'�?������ ���8@��m���|�BL���Ts�O���1����T+�!b��6>��b.,4�e�It���?,ǿ8 f|�Fl|jA`�P��ߚ���6�<��΋�,Ii}��c�����O�XK�s���!�N}}	.3T	��|�U��[�V�U�`Om-0c��.��d�Q�91��<v^k�%=V�+_��
�v�@:�ʧ8o�Y�э�;QGΩ�K2yV�'5��aߝ;$&!�U��gQ��(�*q�$��څx�3gs���,�:$�)�����q<�W%ʓ�N��?���p��oM�Q�g�yz��d�q�+�N�@��8t͙s��Si@Ԣ�,O�l�p�5ր̰$�zi��ڹ!
&{S3����Y��s6���K����ڛ���Xa��!?�{����Yl06��PD|&��R�R"�/=s��j����E�/*FC��@Vo0�$�:
x�?��ڏq�.�c��T��X��C�y,�!�D,�UkfT*���癊��7�.��/��O�M�J�]��B��u+Ϸ�p�{�|���a�|���J�,���x���x#i��"FW��ر���'x6��`��;$���0��@���l��C�g���u�ӂY��VEb
t���%���{��?��j`Bg�B����Kܒ3���|g[��	�ߝ_�y����n'�F�5��E(�y�xt�&���vY>|W
H���L�I�3�2�ȅ�\��LR!C:��!)�8@B�z�Y�ڀ?H�2����:Y)�ȣ�3���OC�F/
��z���1^�B��@h��U��|�C7b�vI�!�����f����?�Έ��_���<Иy���3|n%������m��b�Y'x  �E3׃gk)H�]#�a��T'��ˠ��A�������c�B�nT0��g��D��k���ҹ�<3QI�4о:�T�Ҩ�<�����]};��u ������ ��=�[�ClB7/j��á�#~��|���N�멿'L�o�4�H݉��jK�������f=�oT*���e
8����T�lG����U�vR���u��R�����<*_����gS�IV��	�	�>++2��k���'5�>��@CUUu��2�"kW|�������4�z���gb�щK��1T�BO2�s��z=e�8>��͇�;p��<֒7B��vAҹ�xN��-�{٥�=�=��XC՚Tq�U���CW����l������⨦'��*�hّnSz�A?7�8H�؝�"�@�$E�OҜ ss�3�Է�=*���^�k�gJWV�����Dپ��"�,��j6�M�s��X�a�g��nnd>�~�I�KҴ+m���q�L����>O_����U���K���������֙��5���/sY�H}��`S�C9��
� �ʞq?��_��d���S}c����l\6��<�+J}X ��qo��#�_ �o�O��!'��g$B�Ar��P¡�k���eY�К���EEEeɧ�n1��<���^�߃|@��x&"������ޅ	��e��8�n ����`�DXh+��Pn�F�ʫOC�]R�.o�I���=�TF1��6팘F[�	ba���g��ܟ	r����ꄾԼ�s�� 4=Օ۵o��{
t�~N}Y��ҕ�9�M�NTa/�A����+=��p��TZC�Y*5%�U��]��
$���ŋ�NoY��wa�����'::d�G����� IAģ�.%\�f���D��F�T���!6�$)�>��q�`ۜL��uTK��wW�e{hIh�w��x�Ɇ���xq����Z^�ri�9kkpzo��?�X���3C��
Wӿ�t�F!&�t�d�J�p�/����hV�Y�«�hͨj�UTj��������}^D��C��o ��J5�� Τ;��^vuh�u?D
#x܄/<�j�����#~A��N7b���5���jo �#_���ڭ�!����X8�?c�'8]���hZΆ�P:@�&4�����9X}�ͱ��`��(MOۂG3�?TPxVJ�� �i�|�����9.]�x^����t�G5@�/��ؔ�?W�|c���)x��9_k>s�e�K�E͙��� �𾓸���#��s�-��Hd�4Ia�ޅ�,�sj��^ϤQ��ģ���"�H�3	�$��22�k8���.��d�9ƺ���h ��&�vחu*D�`��h��ҹN��c��a�a��C�n��kr�+k~�'򛍾<�3>Д-�!�� �w�����7nv�y��k�&lOM|rFjq8�ֶ�%T't�Q��n�Z���>mH��xx��~{��5
6�MWs@��R�Q��e.�;)ǭ�O�����\�|k��)u�X潙�{]>7eA�b�y!�S��>��E��N31Х��pu'��s��\%�g�D�,����-')x�״��P��
!�* �l����c쾈\`c�_�D�X�:�T�q�����
���)iv����������%�T�9��?S�årA��^� �����ӧ��V�k��e��8VO��`ˑ;� ���y�Βj���Z2Xj/������:���7��\�ߵ+*�WUW�0HYy��+"+݃�b������f����V��{�h4�����g�䍵�y"s����đH>�d�j������g3+1�ypg��T��y�$���Fy-�h%qee�/����J�����c��a�yG���� 5���.Dc�N{�O_J�\L���8��ND9�1�x� ���H�����'��(�+��/���}���1�ۘھ�P���~�̅�z0h��j�CB{|��="�á������{�� �����R��ѧ��p\	e\�=�IQ�תA��E8���t���h(������M � �|�z�C2�l�ċ��^�Ƅ2[�8y��� ��7['E!��&d�򄇇���HЊ5J2��j0=j�.V����{0г�{�*�;���`L<��ߒ�r�x!��q�}��=����:��즅L�5k�ɒ>.��� [��x7 E{\O��p!�I�����aE�5'ٓ���]�H2zQ
��ܧ�;|�˟��T�^~�3������h�叅3֭�Ė�_h6H:��Q酳��-�w���4�5QM�{��m���=J��Hb�.9����((#ㅃ�<��՛t��2aV!
�0���ߠj�Y�QP҅q(�������;`!0Z�JO%Z�͠��d��p�4�=�+�0kH cU�)$�5K�� Y;�$����>66�><�u��{@=��,a9K!�?��T2�T	��F8g��ȏG����sEqCm����%��-Z���vF�.�MC�Y�)����\Z����Bm�s-�Qn�>.��ߓtT��0�����q0AP�.�F�R���NS}_��u�C�a,��/u����3����:����m�I�*5r{0O��"3����$�����d�lǪnK�x��G�F���|@`��-^���&Z"2�Ni���Ǽ!V�����ɠ��Q�U�����T^l���_=Z��̑�܀b��N�n�D��V!B�����j�q q:��e3�A�X��O�0���q��p)���vou&��c�+o����-�+Y���P�5���?T®I���zD����Pe=u�*�k��F�ڻ���j3���nD#0� $����T���錵��]���JY�o*CX���q{�W��Wut ��Zjjjk7Q�����h	@x-�g�@g�Z0��#�?-i��ȂDƭt����Kl*�el����"�:0��T���<��5Y$zmIVo	���'7X�6m4�l1>ot�p�O''��|�*�뼨{�9��r�x"�ιc��C�b�~W�}�<��P�?|���$�+�uK:��}�)=@2o��I}���#l/�X庭h~�Gm!����")���[����n{̐��m���{�#C�q8WWמ�<�L<$M�*�[C����G�G�w�i 9@8��c<�̡	d�k ��)(�o �2L�ci��ÿ/�K�"~�6�5�5�)��j�ݑ곱N+q���݆_<�W��]��g��X��h�|c4g��h��ܓ���hE�X��C�� ')m{�䚲s�s�'��x${d�IR��z�E�����K8��/yW=||4�K��[���jw���Zf�ؗ����W����z�U���
����?�ZP����FLڊ7����ݝs �9g��qh~���f�c�@�{o�����>�Vl����ޡq��r�i���52:xي�8��@�}NS�C��当�U���q�1�������#�w��v��� �#ͪ~��#�A�3�',�􂙦�vz����l��]��Z��
������ГÎ�?��m�k�v7r��Rv㵣\R ����r6���5�
u3�7HŜ�>W���V�j�/�qA<�<se�P�X��p�����s���Н3�_;���6׽�&©0,�*o��ٕ�#~ub��<c>#�������3�Sp������%��ypYt���4�WB�{z�4��֋,�J��*��g�s�C���>��R
e侈\􆃸�����o���Дuץ�|Hv��0`h5�y-��M������{y�L"�%!7�h�(��%C!�z���%��5Ae@duHZ�Z��`#���p��1��zW���'o'j����T��\�ɱD>A�
��pp�<2w�@S���*���0A���W�"�� [
�l�6Z��K1f:{�|�6����]��kr�!����6ԇ�x�?��1Ш*g���s�6)Vy�w��$D����ҕ�e�Լ�p�}�f���-���Z����}s����?%�OǱ�q��n��dz힒�o���6�o�����dPP����or�bˉnЉ�M�>= Ͳ������q[`�0�����)���ZP�����H���2��>�Eh���D�����Z˧�B������_y�U`�c�0(��|��pR�n���OS~�")��j�H��F�������� e5�_������IeL�r�g7@j��r&��֒�ߦH�v��O_V�S��sص�SY��o�+���EO]�����*y_�~Ѻ��z/�+o��� L>�
�|��0���ɇ, ��|���C��� F>��|�����ȇ,���|�`�C��� F>��|�����ȇ,���|�`�C��� F>�/�0�k��Wz�����K-v��z/� ° �0,�	|�j60�pz`�A��;0�x��ON�3�&;����mu�ӕ5U��މ�{x{�L�_�5�}�
bSE6�,���1���u�ǷG���v�RX�_R�[5o��2�w}O_X�ې���>�r�"QN���)24S�F�V��0`hX���$�����8��(���9xvE�Y��PSeg����B6P }8�k�$@S�>c��c��e��B����8KE�c��HC��P�Ѩ�F�B�Ǉ�'��V����<�/��P�T�P�_�h���&tG�FI�c;&���~�>pa�{��%TEa3��}ӧ*PՃ�aTz�G�C�s��$�|���SV��AOx3�S�S������ �[�p���$�|Lh�	�ZW��m' �T3��̞�us��/�|�# 2\i`�ke4'�h��'s�y0]�pc�8������ɑ��u�e3��i��/BÂń� �:�B3��?�=�k�uS����X,�B����h�X�����K?xm͟*�}������?�<�,hڸ��d.�2�R�����9Sb�`b�aÕ�A{r�d�_�/�����+@�T^��*j��G@��y�m{.��A٬��ݝ'���Ȇ7�35^���2k�X�Ck'��X��"��<�>���ԩʓ�l߸�F09J�N����5�v����r)�Հ]�*�jΔXG���`�'A��.
�L�������·�)��@/��/���&'}��Ird�,r��r�����F��uA��6�x� �{� 9�m��^��n#@�wr��r�����Qr�E��|�D	��g�ǻ� ?�m������F��y� ?����7��Kr����x� ǻ� 9��r����=� ǻ_ @�wr����x� ǻ� 9��r����=� ǻ_ @�wr����x� ǻ� 9��r����=��R�`��G�yG� ?�k��u���F��6�xϢ��n#��w~�g��x� �{-@�wr����=� ǻ� 9�m�y�3��4'r��4޵	E�1$;U"����$�ד�j�ZA/^���o�"A���0Bg�d�f�9?;�i%����L�y���Ĉ������0��ĐC4�Z�=�ƚ����&zR��i���˳^��ʉƢ���(�q� C�7o���y�[������Ҿ����Gm�H9�@��p@�La��0�*�����}6��̅z�����%^Ê89��XCCC<�7 �If�y����yysN�]�󽆙�Y~�6�<�l��rv ��#��²rriJ�BN˟��Z�g�z�˗&�u��cҙ�eP�'GG��,�3�աD\k�%�n:@�����W24�=�u/�7ۉ����4��
e����(u��KDH� q�7q���}NgM�<�:�wjkoog�xxv����"T)m�����~��l���� ��������i0�4:����	f���o�</.�nt�AN=���')K��`���8�"����\�O:��6���0ip�i|�h�h+��$J����i��f�ϱ���Z&�>i����y�*�FDڛ�[[��M;>��?B� �&���H(> �B�Y�M�����}I&i���3�8~���f�g&�$�x3М�aVCƈ4:��˥�@��:�	(����UV�I<�y�/ 
���Y81af3:|�,cH�u����d�p�)"��^�\�d�=CK[���ɩ��JXO�0����f��4���|�)���4h�z�$�5[e��$�/I,��c��ߔ�u'��������Zc<�K��>�(���7�����l�&�Eq---KD!�L֛E#Q�x~��h	�+) n��xBx��%�87��d�/�z���F��f�����mw�q�8�8m�����]�{���6�M�D82+�3�H���"%�%e�ˡ���)����q�"}8w^g�t2-z��wVJ�����T��))?��6���0����8�,н��ˊ���+���I"�72#f�����r�E�91��tGg��{qn��s�ٗ�x���VH�,�Y�rq)��*�0y� �˿~�׮����WV�ͯ�Jn��c�/L�^�������򐾐)�t]V
�y�����ZB��_���2��1��x�>��];
O2�˅�>��TUgY����[�}��C��EJ�EEC3�����LU�������8V�}��p�5I���;*?>�X�{�7gjc+�*�{�!Htu�(����i�$ �`SEt�����D�qrV�:ud�Ny	%խ��e�u7�Y~gg��㬏��EK|M��eo&����O�O�CÇ'��27�4�(����x��;��Gg^�Q�E��5����w0��©�h��G�N�L����;I��-��#�漳���ģ��Zn{-��3׷�<6yY�/�'�����y���m�ݸ"_��܄�FO�m��7{�v�r�p�՗����"�!_�3Q���
�/r��������+��Bñ1:��FN�,��x(.�%.���������?ė&�O�Hh�+2���&yf�<!*�j�n�_h���KN���j,J>4~G��u�"۩�Q ��*�P�U��^/?я��x	�_�/�A�����u�U8�|�~���]9�bb�}�X�m��W�޿�BsS_��w\��m��T��5�ְ� (�A~|A�(v��c�o)VL(ǭ�� ʵof_'��N�ۖ�$��y�j�&x�H���m6� ظ͑=-35���zS8�� ,Y�_-��z�lY����g�D��1�p�����K���ɖ@6 ��EP�M�z0Q2dl�=��Ǔ	o�dR߾+��u�E�8�{�qұ�?�x�/:�>mB��]�ȳ�o�v�e6�`���^î���^:Ɗ� �V��/^�g��a�+:��㰙?��ְ
'�4�a��v���ʿ|K��`%�O�@H߫B�|�xP�CX.��,U-��d��b�D�+cl���7S	�Rɏ/(�!�4��\iǄt�)�E��l�݀�l�2�A����Ŋ�ǰ�
���F[�ڝ�јZ�e��@�2Ch��,<nR�$��2|<"��L�G��
�?�Jd��`��n&�A���c {���fvp�Kx�'�
�K�g�~+��1ko7�9�NTɕx11��r��P,��8�s2\}V䒳s����rİWdV���Xfj1tA�]x�ˠF�gفd78U�I�7A��n���}t.}�j���gn3�c��+H�{[W���$�#�1�'�Ԙ���~i��߶N{E`��gS��뒭�,�~|�Z_�dzcVf@��)�ۛ�^H��/l������P�{H�����첛��4��h	�Gge����j��O�2�Q�W�""Q]�k�������z��1�տ�v��W�t�}�C��I���j�W.$�<U��u���@�%�qg�.{��;��|
f�)�ͯ��B�F������Q6Sd�`��AUOaG�t>�T�����,�{���ؘ���(bE=n;f����(!��>��j��j��fB�{x��
3����Mj2�8#�8i����2��e4�"�tǜ=c�̀uxbIE���n��0ޑ����>��{=�eR� y߹O� [����uw����������P`�:N��~k�S�����۶���%2����
.�i���aAq��ڿ�@N��Ά�6�s���3K���=�ϘRh�Ҡ�AB.���Z�xK�m��ا��&&��)k\/���H������P��xb	Uĕ}��(}Ƿ�%��u���@ p�n��m��R~��0q7��ߍ��ƞl��";s ~ODz���O��75�.T�PA�/�ٺ�M#���6~ �V~����<�(]���?��QAG��|ߨ��Zj�]S�bH�ֆŵ82�c��������ge����}p�i='��T���η����i�_��%�Cy����Y��C��^�����K�_�T1g�ֵ�ÿp�X��3���(�(@��R���j�w��D�����)���/�Ѻ�V$�t�S�`�i�bsyf�a��ң��%B'E��g��#��V3��E�_�B�x������W���_OU`�[�Rp�+�˧�ī� |�>0*��S^2����W���M�q~#k�El_��-i��M���6�.�Z��������Ey���LW*��Ab��IPf9\KL|���	B ��<Cޏ������@�TڦjGy���K���}�S�ۜ���ͅ����)tĕ�sS�u�i�Y ��sS�f'9X��|��TX`�Q�1s�^�k޹���7�52�
��"�6?['�T.�!пE5�/y�N�_�NP�������w߯kx�E�����[U�Upv��� ���^�Y��N�~Ne�iD�C��(Y�᧸���8���:ab��V&_]e�"�tf�B`��=#5�N���lvP>���6���ݞײ��o��Q�����n�M�&��'U9����I�`�����~��� �;_��׶���~��l晦�Z�D�2g���;�2$�)z���U��:@#uz�5�h��)`�/��6v�w���b��B�Qχn���P�wr����vB�������V��v)�n��k�u6���
�Q�)��{D�����E9@6sί���yc�,���g�2�'��0�;�V�[�
;Mw=Co��΅�j���T��V^���˹�f)u^1�"����S]qP���ΌY�r������9�V	��	���b��ؘ�
EO�� g���f�ϯ���v�#��_�-�@E�}����(����r����cX}�Cs0��W2��}��2`�����w'@ӸO|��<ߓ����D�r�]�s�s���v�XLr�n�m�E����(��5բ�Tj��HrII�lIdB��(�.��PӔt�f&�I5�{�?s��������{�8�&����|ݷHtF��3�jbB�Lv�����hcЉ/ա/�Nv�4�u�x��_������,���aR����m�h��������F��qi���I���~��W�s��n.;eu�t����.��b�n]9r[5�.�V����j�����k�����+�+��j�����iM���g9&���-��7ؽ�����%����9���Mx/;c=;�]bo�&$<V���P�GKQx^���]*�v0eu������bA�b��>��������
h�D���+��A��QYl�A*e�UP=?uww[i��f�P)b�Kӏ�;��a+(�����hem]0?��I1����{�$��tG��韏w��U)a�~)��?d���H��8�j�b��%��qƢ�L��ՙ���WY��3x)��A�k��a����Lvo����xD�Pʐ.�l�1�);_f����A	A�'�)t�lY�c�G��D���&�����YǇ:����Q�L�4�q5��տ것4�OgR��~{&lJ���y#�/�]��Nj"&a߳��H}���A��'r����Z��יC��Uo;gT�a��Un-��a���� �w��@��Q��x�c�&�Leg�TJ����cXܼ�Q?�Csm���_( �¸���
_Z7��s�։��&��)�82�zq��qE2p�=����H�_�:��C�����o�Y|H�%��*���n������3I�N�6��x?7�(�8�ʻ��	��2��<���b����G��&�'y�K_-���~�i��بR�Ԭyy�sj#�.+��'�����L�ȵ��p[%L32�匾���dUgL}ͣ	 ��I"��C��¸��G��P������S���dgf��`��[@���2�J�P��e�f�d7ned���������W���T�����c���:���b�y��)<�w��%p��:���5o�>0N�_-��H��,��|�<6[����D�ρ_0�J�B^����r��ei����B"�B�B�}lm2�r����@���mp?_Ĥl���
1���7�ns���k��eT���Zs�$l�vw�_rz�"��\��5���!��qL�����f��-3VM�(��W~d���	7i�N�v:E�X�������DL�y�꿃���۪o�.�<�JD���u����V3��N���	1*#�D�A�{�Fe����Ԁ&��ahpV[QD��&E+�p8��'��O!dd��sn(Wdyu��y%,l�7�8� ��/}��<x-���G�M���- r6��\+��qo�NId*�Q���������	����c��sm��^di�Sq��ؚ����bIK�V�i�ơ�/H�C;>������v:�~#�����\�t�����e����w��Â+ao0{�Ib�<��^�f��Y�ĶL 5}4���jH���K�F�xu.�X����������!�/�!-.�+��&�-T
e�4����?��y��+���#��qp�j���+Ǥzk�ӿ���J�͂�Am�V��^ ��7���	��$��-��J?6N��#���0x@c*����Dy����<Q��L�������.�p�[L`�yMc�4��9��50�Q��ƀDK��mT��h����@{&�����õ�\������޾��#�zϹ�{U���%���Ɛ�}0a%�"����&زoc)�ܨ�i�O�ɿ��q����%Y�
�]rml�s����F#��;cFҔy���z.��c�v����}ز��FC��ի�{��<\�՞*'�"�b3�R^<�;,�&lG,[�y�A"�yh�ùj�s�@��h�D%O�O�r�d<j9 �|���d{��Nv˗���y"�<8�~�[b���g *�x�]�Y��qf��bB�CW�eőc����j��[�"dL�'�>���.�Q�3ףO���ra��K��s+]y>�.i}���u*�J��~wͺ��ٿ��8ް�R�Ɲ�.�����P�fE�:Ѻiuf��scZ��aRw�񽇶,1���S*6��g��c+X��F[+��_���Q���Mio�E��7��d2�7�+L�%]
�Hjll,�}�y�^��&��8K���c⫖��+�K'�ص����WDQ��m֗�c��VC !R��ʈَUi�q���AY���04h�%{T�/*�'�`o0�j�5�~�I�d�1J��nF�GRB� �����[�w��6&�6��RrR�𐊦�hA���7�]م/�t5��QZ��-:�p����]���xV�}��������ݓu��:a�+�Sm��ߓ�m���K϶�'m�`|p#M+~�����퓾6�N=�!�{������T`��_���z ��/�X������1{��^`�����4���O�ٜ��e`@���]�&�di_=�o,an~v<q~+8a%��+� �fm_�L�VH�~ݒ|:=�+�C�!<Xf|}��H�		r�U�ǚaR��7�؏�	I�W�ۛ�K�>^J��+�a�$ѳ��$�UxR�"c��\�^ͅ��Y
���$̥�!����Oo���0������w��ϖz�f\��������e����q^����\|_�՜?�׿��6��@P�|�q��%�����%�8�c 89�dl|�L�Z��iǇ�5�_yq�"c(h�"r���轫e�3t�I>�U-=��m�T	�FC_4��%�}o�ĺK�pѺ<9��,��c�o��%#f�ƌF�w��V��w$���=��~�DF+O��GX;�MD��<S��-�㟫SuHV�
Z ���Fmg/�e�n[
����	�c��4YE�y�\&�j�)8�8���+!UUm��\ͅ㽝���![�~�y�WO�����c�$^\&�cO����p6Lز�qOu���l�`hW�t�	�r D-j�5��������C�z-/���;O[V%�ʼ�1�V%�����5��>�r�ډ��ɗ��_�4�A������ ��q��L+��΄�,b��3�Lz��<�������C���_B�MҐ�q'Y,��yW�<u
�bA���A�i�p*�)V����=i��^nF�N�t�3��3\�4]�]����I��^#�Q�m%��V2��}�.`GԸ�j	^b��t�ҏ�웟��l���t����5X��^`7,��M����Ϻ�NSU[�1v3y���7�����,�Bio�=Y,3�Rv���"N/�/qFOI��nW���q���a@�B?|s�d@�Ɖ�߸M��ʓ�]𕅧�,����0H�4���R�����$��aMH4��T@4�҉%Z�⼱�h��{{R;���S�_z�V�q��g3,L��u�x�k�Aֽ�����#���&��E;�9e�b3�:D��!���5�h5K4�b�X�u�ٵ^g�iQ�:��
��ž�$G�ubIb^�|J�m( ��+����Cٲ�r·�f�����oc����!^^%+��f1��Z�{�-S/�����/�!�����M���GU*4`@<���b����2���y���c3|����l��)){�I4�X�IX���Ջp��"��Q:��/��Y�c��o�1��yu����>���B�[ø"��o������dMV'n\� o��k��V����%�f��?����������
�����i��v*2���?��q���L'�B[�QkvA��_���^S����;)t^T��W[y�z��ώt��@9Aeff~u˙@$�A1qAԏ��n�������+$��#��ǹ:���X�Vy���^ۿH�$�E!���k�վ�'	d��9n(�W�S珜��_Pd	~l�:��>9����EV�B#d�3Q��O���H�)k�^E��}���g�4���iZ	pQ���Oh��((��D�����K�Lڂ��|��1�1��M�*g SϮM-xﺳ��>�s����=p�(oZ'�����[~�2��2�h�kۉ��'%u3�_%A�]62����_���:�4ED�c���F({G�����v���?aI�,u�B���]т�з�'2���]�����Ha���4�9w鿓9O�@�����|����~����b�&Q�ˍ-�B=ɿf�5iza;#'y5#�lW�^G�c5���agе��S�L��`4��,Z�s�/�=Y��{ׯlDYѪ!��M
�o0i����wi���p=�:6�!�sw���	�;�˵w�TgL�H�b�'S��R��U�~�H/��S�4V�9
�����#�ɞHiq`6d�c��_�m�nA�0p��a>������Ϯ+r�p�-G���{B{3쓧�+�Wb�4��j�5�}k���ÆoV4�-x���R@ʶ��j<�H,��)��K��������4o+Ov�کT�W���,����\�1�H�=E�V�MZ��7��q>�ҟ?���'u���iA�}D")�(،%^¬VKh�b6�ʧ����R�b�Z�P*�A5�-�����_�-��g�@msh��D�d�g�z�M���g�o�Ŏ� ײ�^��مֳRv�����0��޻�c�[\i��1�ߡV?�w��X�R^߭�6�M�w*Ϙ����M�dlHE��w~C�>2�3����\�f��m	����l�7,�`W�Mh�c\K;s�r/����`%R�> _Ew��Z1�5 ���n��l�p�F������+��
�b�[NK��+�3��ە�M Wb"���M Z��dB��@��]4��ŗ2,�=)?G�&��#T����T����щU�w�8&`��O��J�o�ȧ'���aƿя��d�yo�Z�r�&l/Pxv(C�҇i$`�^�"RN����)�٤���n��1����e�
OpZt��K�|CY�[(������A����W>�L����z� n2Bo i^M{E��<ɷ��
I��5�^���
��������C?_�Y'N�%���_u��#�s���谱D�T�d��p)�4��b��y�r^���Bc��*4�[����ys�ل9!�*�$rh�o�3����E�`^D;�`z#�ͧ��F=XD�8��/�(."����֒ b�_P�cLm��pme���yD�7���L`�vjA��������%E��(�@�C$���q�Q�fy͘l_�>����j�%伌|Ϥ<�d8:��T�!g� bA�6�[;�A� 0��,+"�!�9�m3�IЖs:M�IKc:rz�����!��L�t�����5�Q�[F�F9.�	�{��&ԊH�JI
�a`��{��Cu8[�RP�]��8[ف���F� x�
�hB�7����#M��oZ.��^|U"�qV��$ �F/X��7�_������P\���(��Sa�]�t��0�?샵�f)6w>��T��7�:�
��g+�h6Y>F�UR��)x$>z1Zml�T���af%J�/4�JB,�?|�I�@�.�6�-����?�˲#��N^}l�-eLɷ���ඩ�m��oK}�d�����i�T����!9�3�^���aY0��%���s��53�~/�?W>�iU<s��n���Ʃ<��5wz_e7����(���Sbv��ל�Kc�!�g�pb;�������~��p��Z�i��5H~�]l���ψ�:�B�>|��"+��1jc��W���\���.�xH .����Ue�7��������$�-�r}���cc�G�h�8�vEE/��Xqc`~ȟ��"�xz"�a<ϓ ����{�SP�4��V8B>�33>��x. e���峪�̠���X�&×G��we황9N*e2L� ��̇��f$cm$v=�q�u?�*^�h�XqD��ݦ��".�1xAxk��1��xLq�j7��9��v�������~�� 5��z}�I��[��4Zɨ�Ȑ�w-��#�eم��߽0ި<%��d��<$�k�*��_��Z��o���'�������,�߳����aK�.7��U���(�A�t� ��f䝘�00�|<$d²
�dY�:���`GҔ+�pË�7a�`�&�/-�,q�>{����,�B�°�.���:��x;�  zO���N!��*�ӜFk�%��~4��ݱc�����2��^-)�//h�/�6�ٍ�q�+��-��;%�#��1��w&/CK����BZհFk@�bYFF#.�J�W6%y��=��1	,z���H��������Ԉ�C���%�87��p#� ��n�����(I}���m�ݩ��Ldb˷��N�t}Տ���,����0��8V~�Qf`�ʱ���b���� �1eb��ͫ�x�;�^^��n"dT5���^�6(���+_G�|�ǒ/���x�pϩ�=��T�U�Ć �� :�4�h�3F�-c,�{����&��B&��4?E�z�Ec��Xp�W��D�
O�ǟ�$�&�_��ȟ�܇�<a�P���dD��F�U�T��{[�n톹�8�����0D;Ҍ`��pA;�1CC4|�B�������K���I�g�)�TDuG��)y�MV�R,��n����w���c�K� �3��Ow�)X�NQ�z�gX�/ X�V<�S��|����8_q��a�,9��`)Ԣ�������D��M�>����3gZE�/���ţ�c
��ѯi�mp� ���ބ�;!O�{.�S�z9�Rh �q <@�N��*���U���4����H����PƑ'S�`�&��-*j���m |R�~|2*Ὢj��t�(�v����{G�����h)�ӓO�$@��*c���r�r�[ΐ�wD�
Ԕw�X�\���p`7��J��}<��1�8;�X�WҘ��'�ܔ2/�R�vvva0�VB92��ʚ����u�	D���`���2���e��_3:����$Ӝ�=Ch)��)!�(��@af�YK�W�!R��H�E'''��T�n�(j1G��0��^:�e�Y����Q9Ɠ @�0��yh��4�FK��Ǽ�>cd��li�E�/����|��$�/�^�H�X^s���S��M�	j�K�B�C=���*g�QMd�K�l�i�I�0���F��/bT�"���N5A��h����1�
��	Ӟ�]��IX�������Y)����y����^�Ղ���c��ݧ��{@!�!̥�`N�ϱ��=1���n�#(y`�-c=�&�� <v��V�ޗ@�7��������4����_�ɏ���ߘ��P$pl�:|c��j����Z��
޻�fA �f��� �z��ZiS��1iS���#�U�|�[�- ���)ɶп?���`)j�����'|�o�On��χ�;/��4�(�����ϸ��}�P�}�9H���2cl�Y����Iw~[�cɊ:��9v��[�wJ2��Ŋs�|q���1EEE3�&�[����b�*���<��L��D�O�>�@��<��I6^II2��B��S|$�	�~��w�1-��9n�����}Z[� ��tTY���s �'��ҢGV�]j��R2���w#���A0�< �U6
��ɰYR�`	�:-{xw��G��A���0���C��v#K�"��"b�Ƃ��D�ٶ�+�ޯ���-�'\���I~G!Zy���W��$�3�4��x�����a��[�Y4�vȍ����{����,��_��=+�4$b+������b�Y�'��vf���/����.���c���8�o4�6~u���4�8D]$"��)���Qrͪ�K��6���&g>^ʞRZ���7�Ma���B�8|Y*`�<��^q�!/.�"�=��=�)�)�B
U%=f�^�!"L�Ω�I��%�:^H ��/L��,MٸďH�j&����a�x۔��-{ش�I�������@6ƌPh�K�|���PJ���{%���u�`8�
�!��B�A5�Ꭱ����h(	��y�&�����y����ݺ�(U�=qJ:�=�':cͷSe�=ݓq����@����o���$b��Da���h�മn���u��h�H2 Nٳ+f�#3��,J�y��}n���բ��V)I�����ǒ�ߑw_���;V�{�=�^�d��Rֆ��c-^���bwi��%��G	q?ifo�f�|�xyPR���.�����8��GRuWn��������9�%9#C?ncqEC�����J�l��ټ#��T|�$Ԛ��V3���DB"+�NVtV7��㾐eu͛/�(�dd���@�t��N��N��Xmz/ٍ���׶�&��a�qY����2o&��G���Ӳ~�4K8mꮣ�T텬%owԒi�rl�C�$�c������M��c�ZA�U
+���by�Eb� �8,��Vx��WB?2r�p_���P�ٷ��Kyx�kR�RZVz�m8UMG,ʊk3��ˈڌ��h�,�k�u�V#��`2��x����ـ4[�1���0����>ֵ{?�X��C��R�=�v^D�!����Cz�%lկ����Q'{�ޙ΅����[�!�c��u��sj
[�f�)q}���}�\M7��P*��ju"q�����u���g���7�=��b�������qN��_��v!~ZR8�e�k�o(�mh0�4�p_��rX��8o58��a(I�vS�2��,�ս�g�a%'w"��
3�]�}��Y�s��K�]�?�N�ב���s]�(�F�n�Cr�0$ˊ�iqun>�JsCY0��H%T9"司�\�3
���Cz��vX+������s��"���D�x�>ׄC�&��߿*j��R.���e)�D5<���Y!U����^��.��U�s����k�1F_�����oߴ��l\r)����+'U��c�����M�I(yy���0��D&�T��3Lj���3���� ���M}Pt&�N{#��C��0�۵m>���ոP��f�٥�&���|ӆ���@��!7E_g�.�X�p9���z�;5�>��q��nm� �-����&�v�"���4�[wf��+U�����g���v뢦Ï�u��	l�k9�ґk���ӛC~B�`5�2�L&3���r#-W|���:��-CN�̉�H_�&Q��v�A���u�J�WÃ�hn�^*�T�Q8��G�Po���� �É?5����I�)�_=s�N�J=�N��jng�T8���
5P���.A�s�2%%`��p,��t[��.���?q�����VQ* �����=}D�c�,������-�g�#A�]�^:����<�9�p�eBR�Q�塡!�ԡ�MSP����B��8!�*�3-��e�CF1@s.b��ƴʛ0��ψBɃ�:S'��R�\���d	|��m��|!T`������k>�hI�E�\a���;�8_Z�C�Ppv�c��آ�R�6�Mu���������ʧG�P9�Z 25~����$Wa32�k;��1L6e���K5�Π�~W
K=^��Lnm���mk4i���ǵ�{�}��	!w��1�굾���d�`�5��*�z�����6B*��w���?����$�W]���`өȫ�sZ$2��۳*$��*��9[^�3�PA���m�/�����0V�١�������(�=�����H��e��(�=�x~'��M�n焘2�_�{nP�Nª8hIvc��������~߃�`����� 8���қ�e]ߴ^V�Gf���q�($��^e����S�&V��utoH������D��T��Y77mz����ݭ��{��ܞ�P]���w���!�t��0O���-G����#6��R���OmmK�s��~:�x�F�;��OS�:Ҹ}N\������{�cV
<�n^�Hо�jy(n��\�<o�k����p �M���$�S�����%7A�UA��?��i���{깅	(���~|.ԁW#GE���y�>n��5;��4��K4䢼v�P˘�m�����dv�Pi�$k3���YđA�!Π�j���آ>�e���Pf��Y��_%7�J� f�� �-g(�{�cu"j��������C��k{�,cy���n��sG%�F��T�M�73�Z��"ċ�(7"�����?�����>5��g��e�_m��@��\��68Gc����i��6���r����[��g�7NG	d��)u���X�xU�(�l�|�n��p����uJL��DR���̔� �>�?�yK^(�b/7�nr�<�3�]j��<LNNb�۬[U&#4���'�S�O�_�9�R�a��y� ���^ؚ��{�T�?.MUo�_�8��B-��](��oH���lݭq�։���1���V���M�@)ű,p뀠�vP �T)-�m�r`���Ȱ4e������:iB���nBE�c��[�Аi�&8w�k0�Fx���R(�rJ4Q�Ŵ�W���u�%�^^�r�}�����ڡ�_F%���$Az�C��dC�H$��ǻ��� ~��\�V-���G��xA�4�ڨ�ګ���e�Fl���_k1����G���W��%�
ZB�sW�z��^��g�Zlbw�	Y;�y�P�4���P�׍��.�g	��(�v<��J'�[���\�ѭ�V�%�G+M��Y2|�B�ת-�+�8����Ft���:�L�+�Óհ��Kr�7<z���x/"�(E~{��-�ם|D�z�K�P�*�{�Y}�z�UoXH����[��J)��O�N��RB�,{�/`���Cb~�tVX��`|F��\r���R��70��A�a"��K�aPt���v �ߛ�2)��Đo_�GK��n��>��]۬^]��(UL���`�䷚ۅS?i/�F),/�<#X� -����%H��-���(���<�@_��~�&�CH�ң�-ZX�ΐz�#��ot�ڬ}cJ�]�"���f_��}a�
�|Y�c$Y���h}�cog���+PR޹/�.
(o�
��XH����O�>�H�͟��h�jS��lmJ������`�> M��;`\�`!?���g�8�,Џ ��#޴G�w�J����̏�H���3�6XB�ؓ���q���Yj����h�_�����h
���29l�A3`�]�օH���Z��se�'?�=`���Ϭ�Z����[@�������W����?�vD���F	Y�\��7�<����;'���m`A�oCL������W�j	�2T`^��&Ɓg i~_�&�F��Ί���3aR�T@�M��K>���,hu��F'���� 𷒦���i�7___��i��]�/o�p�������3�~�:ckk��њ���ð7�x���3��%|I[�O�\�tL�|*�7��R�{8�z���	��Z8�qUj��{Ξ�8'��k������g6d�
�;L����?��!����u(m\��Q��Õ���)��/j:́H��{��Fee�5�x���+����:�z�E��o��`���yα�*�bt@K����:ʤ�ݏ�D��R��:�]1p%+������Lھ�X�ֺ~�!�HnG��~u��_�R� ����j*�܅d r!�ˮS
"fv�w��[�R��ez������c�9�b���6z�^�V��y�� [�ޱ������'3j��������f�}�����G�36co�1��pw(m+0,]��9Z[%ɧo�B��)�AP ���,�ڛ��g �T���҈RG� �JS@r����^�<	�C�AU�Ѡ�!���ʸ�TT	�F�t߅�$YZҬF!�y���zq�7�H*I��p�߷��-I�����S��=JUw���6��pml\����B�h�0���֡�X[��^e�9t���	2:�{k,{HE�����g����5�uϮP4�2�/8����]12��9��Y�㩉�t��r9��`������22��f��i�Y��a�1�2�S�3#�i�Q�\%	�n�����o(�)ة\��o���^\�*JR9���}`�wA3H�Z�J����J�����g���]y%��I&���L؏�=���ި�0��E��o'�|�A��8Z�av'��/r�S
�:7��Kme��bo�;�	�p'R]�����?I�h��B�nUU�T*4ak�M!A�z��a�|Q�$_��e'�<I4�!�ץ��"���i����Q#���Z=��n�ē�Yu]�l�G?�1�k��j��蕌�bSy;	�=]v@�îS\����׬a�}v�j���W�K����o,2]�t�p1j�X�%��ϵ�I�y�*�m��F�kM�:#L��[�|�,6�0M+����3��(�牫n�-ɡ�-�=t����m5�59����l�ݿ��Z��o~~>���~p?&����wZ�dD�K����\�"���s�.aVCU�s��P&���l���V�d��9�� "�S�srr�C,Y�� �v=�h����=u���Z�[|P�~?	M���bT+�w��������YŒo�R_� 9�1L2��e&��Ϟ9�]
��Q���ߖ���P��m�ď���7�Vn�h�W��IX�R�R�Q�4]ǲ�[e�"c
�oq˝�L#Y��g]^�f���k�a_fbO���,�	�����a��ۖI�A�y'������nlI��� ��d7�3oR��L�q��$���Jy�qŨe���үBS���m��8���؎c�7�:�D'o��a�G�̷��J�6]�]1�T�������e��
�0�Y�D�7Q�*��j���K���7��]�A�n��	Э����s� }��|!���S�UJ�2��ޑ�g�R�P`�x�U�NJc�)��Ⱥ�w�Qb��}���yv@1�6O�?��-��U��Vy^3������h?�F/T�+�-�A�(Cݵ�5kr�=����;�-4��5��D�-ѫ�v5i�
o��ñw,�H�kA��v^�Պ���1��ə���Ǒ钦����8v�E�����	Z���t|��7\k�E�.Ҏg��o����k�~vej`��U �X�=��L����_ �XC��꿺��R�R#�wh�U'�+5��Bi4n�.��3�+���oJ��q8,���n^c.���t�P�E�F���᳹Ѳxg-����~x���fbn.f��wvio\Z���%��m�@���,�A�1����{]�C�v`���5� 07�����3��c�K�h���x����+��kف�~fO�9�����x?!ҕ�+۽h�I���v�������jl�h�8������֣���A%3�3#5��Hu�t��ԍ_g�7[[�!zW9����+�n{���i�sԓ����h��$���@�_��=���'U{�+�2����QV�f��e����7�Ji#_�}U�?���Dz�j�� eつ�����) ��g�����T;�K��c����3�aV���p\��1������Eht��,<r.�=!�C3��32(;LA�VK�����
P���r{;��֦nA.I �+�Ʒ!fXj@R�z�jmA�u�
���ڛc�Ih�W%���4��hۑ���P,j�����l�䁕0�b�Ko����O�f���+Т��G��RcW���/뻵�FĦ�6t����9�GR?�_��1D�R��sz�o}������␥�3�_r���fd���\�Z��'>Ӵ7~��1�s��z����&~��
.nf�IG��*W�`�� #ʌ��r�N׳��xԊ������ t�eC����=�,��'�W"�oLU�K'������բ),`E���J4�I+8,�yuŷG9YYb�r
�r�Kں�R�����\˕��],�_�w��Y�N|�����pu�G�v���<c�T�Wb������w�(��Cc���oN� $�����}����gצ"���q�`����o<M=2o��"s�^�	�����;&�k����z���z��"/r?�:�8��x�������+V��nx�ՠ��?�����_��٥�^��:X����(�ڃ���_�����|"����B������K)��wơ�mC|}%�,Y�ɍvX�s��!�-�Ry���n?y��^�-���K`��}����ϰ.g������;���L@��ڗHB���:��CB�O<�z���N��^�]^����4;.��`Ņ"k=Rl=�)=¿t��A���i�����E�����:{0�(�Qż�]&��(q/.O��G..g#�O���vbߔ~����ĭ�͈֪���5Hn�xRW�TY��q��?�����IBu��N��ܚ7tSO�چ��W�KKɏ35��������ΡK�Ux�
�
�v:�N�Q�%�"��-l �2f�[�WέO�.��e{���fM���]�����Y�t��[c��Yulc��ZZ��0�+X��֝?��u�v�Q�v�ơ��K n,g�2�Y�#pH�S���-K�G��dr	.�{����Yd�[N�2?�U��o�n���I�e� �n�[��1�0��vSv>G͛�E��X�AWB9�g�O�%^1��n����sN��v֦�GQmNً��j��E�C���z��/=���FŁ�7 K�������JEI�~4X|�GY�l�b��ͶQ�L��������욠
�;�PRے���j[`ŇA��w[�~+HzD�D��ˤ�Eɟ����d���peY$0�#N�xr#}����5;�Wݞ���R�ɘ+u��Ř����L)�|% S>@�dv����4(�mz�e�!�Mb�����\�z�O�4طg��}y@�E>Y%�{?6 ��9��X��(��o~�rUms�;�^hhtY;_,�]1)�J�ɒoO�%O�u`���7f���@����տp�49쭣Q}��MJ�ޫP���U��#3���0�m[�S8T���5`08-x365��a��.�뒜��3 ��)$�jqsr1Ofn2�so&��c�l���5Wb�v� R׈6�|�_�TVܵ��(��Vy|�3�����:�if��&��}%t��u�5W{����X���i���;Hн*���7��b2�N��LM���
�$��ۻ���|v/���}=;=h�d# {�<��]��-�!ˍ�E��Ǖ��mM[�y��W��Ꮢ|F�����X���O5Q'@�M�4��U�Q!�M����:�FV{[��-��az�'��Z�8ŋ��	��\�8T�	j��d~�	��.3��K�ښ[��_= ��������kB�~�[��=kb����pf�R�b��%��wJ�#�4�#���	+<���C��*_�-R*L�p����㶫��2p"󈵵��<�\2Z9�?������\|�Ws�C9��YZ!	���Vhf���H�8GaaJ�]�V�'���~A������A8+��E�R�{+������6e�G�?'�A-+@�J4��TF|lҦ�Xok��þ,uG����y(�K"�߆��X�9i�D_o�3�W?`r��ea%���ϛu�25O����S�î6d�e#�����$�a��/s���v���z/�N�#��t/��Ο(C��NM�0���21pa^xa�Ԓ�|I��{�[,{�7{���tj*��9z�|4c߬Y.�Q�j�TI|����=YK�.7�⋵�]t�j�Ûx/<�-��m�>G��T���߻~`���p.��4{�T�\t#��<0���l���֖\i��[�6�#|�I�NwX�5�jC�u�p��U~赔��PH5�ݿ ��C�~t+��A����Я��dߌ�m��/�1x����-ŵ;�S�45�8� R������{4�,��73��r ~u"�����7�ё#{�����A+����t�5�+su�x
��T���)��j��_���FZ9@��;��I���$~���k����+HA+�U��-D.<�al��)Б�hU���97��V� k~p�E���CHNt�{XB�B�z����;�XS4���t���t��[�U�Q���6��t�SV]wr�vz_���C�Ǡ�´>��D�!oH�6�hW���v*�!�!{[�㽝����-��Ƴ.*��CÀ�{D�-�l��)��/��7��	�����f�

�z.o�Y免p]�aR���lmڏ䬈~�c����/��n?��BPʟa9�4������Jok8z�����J�o¡��sޮ�+/@V�p��`����ѻ��Q
r�b���Q["�v՞������ܹaU��X����]Y�����@�G��o/c����S�p:k��)�,_�'��=U/���zJ�x�W>sB��m�z���k0щ]%ED�K:�V����6�FI3q��kkVY47�(m���԰]�i�+��U�Ӹէع��#2D�/�w�fA	P�h)�)�1�BOd��������G��q|D>��z���a�t~u%�+�G�j@�Gvzж7L�ജ��v�� �x�J��۔_pH�Wo�`S,vh��y��Um��$�֠�M��c����J��"��<d���S�����3��x�B��Tr�q��n��_:�k�#��lX�T���(𺾅���^>����+���_�W��2:q��?����������%J>�Јi��&dʬSje��>�t�F{�b0F�l��"P�fl^�c�R[�x]�Q�nO�tk�e������L���8��n��@[N""aeN-#'��O��`w�{�yH.蹘�;�h+�h�����i h&��T*3���Ƶ{ᆊ^d5��L���o����Q���Y��Ga	��CMc%��7��h�@��� �S�f��@#�%�:��g͒ތR*���_~���p��[���^NvlFU;��,%�`jr�54��͹K�p	����$��ե��s^Q�' r�:zʥ/krE�0ܩQ��c)�0���������Z��ɗ����B��n&.��
�<n�������"�вs�C͗r�6`>L�^�Z2E��J��@|n��H= D[�E�H�|���E���p?�@m��	����;H����w�#g�Çw����8�h	7-�Y`�m��J+`�_�Z��γ#� gV����zZ9F���`B�=C-�9�C§���Է�80�`��q�:آX��bw�����J�E��a��3�J��_�Q�����4��{W���e

_�P��5��W��!��w��kDr3�d<0%�g�VԞ$ÑB��;�?}�0h�L�|z{p.��K���ۼ���ß���\�p��l�!y�␄zڷ!�!K[#	�.Zzֺ�@AAay8jmړ"9��8��:�fR��h"K�V棬�v�f]��V�$P=�k�;"�e[dRk�!�g���yH����E�f��01�>5�������AJ�/\d	iD$�m�2jq�O<�P�՝{����0�h�{�3�텮еD����������d��\끱{�G�Ê�N��ڂM����E�r�l��!�	�D�`�1�/�䓩���&�����O��G��d�o��0Gѹ���YB��֘�w<���Ո�9&���v�݁V��q��%w�v{�N�N�TN/�@1^&���aB��Z�����S^m�����-#��	k:ZW`W����3��u�y.�ȎPY���݇���N�0�C�!�4�ߠ~�CK�t���fkk^�l�-�JVTI�,k�IUG��N晽۸2���wK�^�qۚ5܋���G�N5�uͨ�JyPʇR�=a ����'���!�nj���g>�Y��[F��ai(����(g���P��<��Ch������O�D��'htd$x9��<�
:.�_�c�U����Aֽav#��*���@T$���5���H�E&�2Z��LW�~�ה����*DZ�~�!��ޢUE�h��~��2���n5IW<S�in�(��=�]�	�\j����h���t��rZ|�՞���e�������НFK�.\WX��e"�<���^����t[r����	1���d�sjB�O�^��ǲ.�1>��)aTϕ����n�$Z%��ۖrJ�L�Q�*G�(��Gݠ���N�"焖�*��9�ps\"���3��W����W5�Q��AK�6@5�EKM���|���U�ݔ��y�:�$��Y]��{���yf�u��%֯�־䌌�� Y軮����� �W�;����+��VCU؄VA����%�BA�"�؞�=�N��;��A���޴� ���a��eB��4$��%��<�-�1h@�[��3�m;ާ�V���M�Kl���v֮�+���\4R������vPK�Q�R��>~�G�=dm_�ӄr��c�B�1LJ�ќc�b S��Dv v��b����M�Ô�{)k}?��P+J�P&��xW��l�Xi8d���:86>��q-��JS�Ι(�˪c֪�ႌb8�i�0�ϟ�fr�7��Ph~�	���ڬk�I��O���eޢ���_��v��6/e��̮vVuB�d-j�k��~�W�Qv[$�B��K]�0~o
SJ��6��D����8%C��4�zm�'5���!�!/8������������n��h��֋�2��q3�^55� �Ov�h��^�f;��ۃ���|A�[�����h[14��Q+z�p�5�f�6�Ė>��U�=xo]uTYK|MB����WwԦ�C�86]�&r�	��B�����Ji,�ۋ�buut3[ն~.�Һ�ӳ��F��q�1��<:<p8���d���A��A-���#�9��ev��Ͷ��n��ȮY("��s���Sϗ�?�p���s_��GL2�!?l�D-�iw���xɆ���`S@`l5�������&h�V���
_�l�f5%Y��fm]8�����	��o8�t�p���t�������<d$H�ٔU�C)�)U���L�Px��UX�Cҫ~#K%fTǌ=�.���d�����������eꤠ������>jdD�:���M��l��_%���8�;Pu�G�����m�xl��)8�¢W�O�;}7��w۳3b
v_���2��һz�CH��[�n&��� `ms�o#���� l��2
�UǶ$z� Uܟ�Jon	)�V�P��7�3f�5�?�d�4�)A�>�^:�Kf��^��b��-x�}��72�׉F�_ۂO�N��w/��z~=�}�
�Y���2�Y���5�P<Ĳ]LJ��+�~���ր���sg�������}�s��^*����	=0ڑ�8\M�Ҏ���	x���!J�ښ:C�Mw~[���������E�aj�����H4�J?Mұ֩�@dR�^����)���s`g
�3�pW����m��6-�Dgx��
7�dv��ނ��PB�l5<�Ւ�WUY[�F���mUa�9�b�I7\�
ve_\t�W�PF�d��>{����u�Ee#ZqR����8�өRj���upx*}�k���ܩ�ܜ#�5��s�l��8_m;\#���� #7�/
_Y��IT٬�8޷��·%r�6Yz��\
-��ҋE h��._q��_=��#RV���7m��뭦hL��N~�T˨�G�h�?@��j�h�-��ĒՁD���cC�r5�8Q������fd`@w� �<ޓ*�ػ{�E�0M�" �Oe���U��=��xf,�qy+o�w���=�V*�N�r�\���(�k��Eݿ�mfz>Q�"����,�����Jh��Ճ_��-�ƾ�$lCW?b��kI��kSmCxc��E�	�@2�(~0�
�W�OZT]����
�e˸/�۸��
�H� Ǳ�p#�HkS��b��og��Z�۩�ߥ�X ��	~�P�@%��t;���n��G���Gw\��S}ت����Y\�t9���+.�yҌ������<_�
M�s�E�.#V{XTw���c�\���7u��b�zނ�mOI55[���̟��8��ve�� �,��r�V s[�#�A�����B�o������bIؼ��,|G�1f65-�,���Q�}�+c��S�x���T&�����H$Pŉ�XP}�9$�DV���9�\;���u����%�Z��ѡw�pi�W�
޵����o�m���П��)�f����J
l�V~����}���qæZ}��g�u&�J�O�В����-�
�xx�|ʉՈ��m,�.���K�Pn����A`�f�,H�^(�g�I�<��6���c\FM&���v�4y/
੭��/C'&a}V�c#J?F����$5{�s�e��@R�\w�P_'��޲6��{�o�`������Y�J�p��.�<�p�{1eee<tr@���,QG��^C���	��{��n�lf������]}�o2}8���z��˧O�;�3�̓�1燎~�+�I������"x�kl��۬S�F����/F/�\�䅎m?ױ��E�ٓ�*��<�6L~�&W<�����!��=�<\py� �^������� L��7 kai����lϩXe^$��Ph�(b�ׂ�@�}�@�gЮ�8�G%f^v��l){`��`�9��ZK-n�'ګ=�h�87� �ò�괪";�;�ǔ���\\S� V����E�%+�l�^��J�}x�ro���dH��f56�����:G�����gv嘹?�n��<�ߓ�sm��E�ցߛJ_ ���L�Xe{/��"	���,����hW===-�l��!�/�ο#����&��v�9���k�����k�l����D�tu�0�0Wh�ңe� m�����=���Cs.��J�t�L|��aa>����CX=�$�}%q�k���繟m�5 ���=����X�hT�@�դ����g�b��z�c�.��`�+a	��~4��´�a��\�B1�1���%� ��uw/�_��9�L�#i��=-�� F(4@@
���'���NH�ˤ�N��r*=���rܗ|�I�	:5�߳h�B�Q�F�yNM}}}.k�>��B�87��S7���|'����ú�����ŋ5�w/.r�wލ�b�'�k�jłȟd����%�0�s�D�z-�2�V!۬�����j
e�O���#��v�d�i��O�&���=%V�_�;B�{�'w�5j���λ�xo���3躄�=�]ռ�x�n�*�n�O��9���'k�v.JΓ�MҺ��/��FP��7.�Ww2
H
�J=&����WUu0w����na�@�n56�q��B�"T�Ooo�䵵���m��jeb�* "A@�VA��`�29!
HCLQ�UDEe�F@���BZ(�"�L"$H ���=�Ы��}��\]�Ū���=<����}N��T�'0
V:&l�-Q�{{�h�%�A�2s�-��/[���-��a<K�9�Xz�S6r�Q:��F�%���B��m6A�FG�1��&B7��s�yܻۭ���Q��E�I�
�m�揭A�ΨB�ˀUڭ�a��	|[瑤,c�決S���m���jN(�tM��Z�U�,%�$G����|�� No�q[Du�)��|��{K�2Nh��؍��I�^�w����6����rD�g�r"JYh�G{K�Z�>!nvC{e_Ӏ}��C]�q�w�9E�G҂�������7��h�i1|�?���'�!����:NT�.b��/�8SG<.��kv"ĸUc�n�����y�F�����H���喤Ԥ@~Ti)�c^����ג���f�u=�b�UVMMM*�z��xJ���P STT=7(J�8ش��(2!>��ȝϷ"1� %�2����t�j�>u���
W!C����5�����#�?��+_���5�2j��A#�@.h�&i r��=�ӲcopݠLS���N��D�)�I1�+?�Q�%�|̓CA�X����26��+�+&��f/)d��<���q��v=�5z.2h������
`�Ӫ�-.���#��5�gfb�LA��/��m���M�l�ŕW�A��Nz��G}R��4���SͲE�Aa���,�;��9xiT�:::��,0��MAv1�ݜt�q��ܹ� 3�F"��2^��he+G�&�:qS�h���k:&�?&P�d����qo�=L��q��2����M����^dY�j9�;(�S*Ȯ�_�Ω��W?.���|��sr�6,��0�v4�S5��n��*��~y}κH�� |j�/@����	,C�jx�K1�����BT[����"���5�ݽ�v�HǄL�p�'���@�F�֌���C�ad��.�"���@����(�Ѻoia��ULjV�t!)l�X����O�8��mR�d1�����=��{#�񖽿���RA΁����� �S0,,uفJ�Z�A�s���3O	<�c8��Q~� yi�X�k%o��zU�|�����H�X^o��]Ȼ�f�L[��1�AQ�z<��m��mK�UA�R�9��������!�����RQX���H��	��o-�^G��ʪ�N��hve�S�&��1�V�b���+є���-1���H|tM��Z��m	��;+|�G�'�P�%|h��5L�Y�l�y� {�?�{A�/�V݀���Ӭ��D�$1O�y}��8fj�%���%1~��N84�'���x�3h}<444o��"���F�<Y²/����۫�c����c�S����%,�VV�J�5��֞h�^���Jx!w'�(�ߖ��`��+� ���g�>Py{,s-�hy"���������5��kB�	1�8fu\f�8��GP�5�^���%]�,Nbs����4� �̩���=+����>gmmݮ ����N}��*^���K�wzG�p۽��I�'��xb�,S�42efl��	<4Y���U�sn�+�Vl0�9���M��%�ds�E�A_�X���	�똨ʘ�3 /���9g�)蒒 /I��z�ftEc+>q�M��Vm��'$27v`�,�z���Dh�ė��bj�u.�L���t�(}/�����D j&l��S�8br2���Dr���g�Ƅ�?9�A�s�r*{?��غ8I+I�*�8�S��w�3� j>����~ޜ�p܇k#~EKf;��]ƪaŨ��k��cnW���#+��O|&	�U�q�D7�
e�^*@zǖ�!ڒ��c�W��2���e ���Cf*�߬XR~�]�|-�~rI��=�f��r����˘����$A$U}>3p �A�yW��Y��Ե#+{V��>G����K)�R#��6�C%���<���:Hk�P+�[T~5�r�kh���S�U�{	I֎��'�[q���o5�05�
�@EE��;P'�C�����V��:'c�p�w�~7��Us5໏tU�s$�n���HܞQ�������T�p�ݎf�y]����XHbe���3�h�V��WB6x*��H_���x@'��;wy�t-&��r��c��ぅ��*�cW�g(�8�0�t��[ɪD�sgu�����-6+�U$�u;B�b�-q�mh�����>=(q���a�A݋�OΗ�� ���޷��@UU��mf%�v7�T5ı9���;�2����_(#��
0o�I���Y��AQ���!1f&�v^2{ot;W��"����$�Ao�Ѡ���OP�ߖ�.N�TsI� ��U���r= Gm���~�bq��T�2��W��?���d�o�e�`S�e�3`�M�����
:zt�C�P40=SԦ7�c��=q���;���Ǳj�`P���y{"%ω�<���@��稠�Q�,��]2f�y˔2떌���X��Km��;X�^R����f�5Pan%֊q��b�l�,�6�lc�i���'H��7�Q{ظ�n�xV�˲^�^��ϥ�>w���n�q�x_�KFl{_ �H@f�(��d����S����2c��-?A^)��mTVQQѓ�Vz}�ĞLh�7��7;�%���Ք�T���d��6j�$>sY�?�,��&'�~��3�Z�������C$���$�Z�����~s�V��.]0�xs�������V�V��hr�Ts����@W�|LmM�i���G�Vygt"��F�8ν��߽w��D�cl���0zV��zk+v,��:�w�˪			Zܟ��.��
�aP��[P�k�UCKt%-}�vX�r���%C�Gw7jF��~�$U�z����m�"Scz"�H0��	?�`vt��c�I>�P"�'�a�&�=��������/7�+�U��҃�ãZ��W9�Y	��[R��'H����� �-#l$��Y��G�l�ˬ"��+<��ܸ�0"A|��(��u�!�XV�=ecCsc���	f�/��'�.� nI��� �N�#�H�y�W)�3���v����Qd~V���+�d!v��鬖������r�4kj��d���cZ0=0�'9�Ǵ�!c�x	lȂ΀톾�bA���w��l ����x���n���
D]���⮯2��̀k���QFf��U������vq����2 �����sP���q�mK�4Qѡ��O�������3�q_u����k��BY���H���o��\Ri��c�׷��w �'Iwrt���i�j_f M����2���?1�=�mNr̢�ҡ��t�`��T�c$�&��[@9���jP�AQ�O�@�X#X�:n؜��a������d�B�wt<n&��QO��ܜ�F�<`D�@?�ٲ"$ކ~*�W��6��E��t(^;3vl���#�V��~�bb�OTgR»@itf]���l���ƞ}����tTNl�Kp������u�D2�e���`��>�5��
6�d�,*~0��)$��M��j���Y��æ���48pnJC�^���q��0�����2tvtgG��\������
LRMRE����^NzQWW�Pe�;h�.���#4��"���N�|Mkǎx�̱~�u��6���F� �y
=�*$b�L��п�]!�`:��A��h͎�7:�I?EM�����NI��G��c������6~��/B�lS)3�=����e_�$~μU�D���l����$�O�	��6!����'�E#)�����TiF���S�:��F�-��X#q65�#
�x�m�NJ��k�� �����~����/���b��(ڑ���f��裯_��I����*Ap=-	�,���җ[R�Q��,)���*�M���-�ؗp����7��� �U&� � �֛�?�i~zǊb�)��CDx�o�x�r�8���}�5����Jʬ4UP���@�Cxz�1Iە!�� �t��?�r1ڷ c�{E�-�eɨJ+߻�ۣ�~�L4XZZ���e2jI�ݷnWϞ�mӋ%Z;�K���1�H�@y�^�����E&p7((h6V�>�x�Y��uWW\�dT�J"Yh5i����� :�L�e��D)y)�Ѩ�������TDNGo@g�W�I\>$��	�D�nrs�ʂ��-�E`��ԁ�sp9=���¦�z�
����g�(Ɲ�����Y�M��(�wg���wY�/���G�|�����VO1Y-�,��6��]���k;��}w�G��=�_|�g��g��>���p��mU�+Ϥ2��D1����߅����8�N5��7�7t�����%�$=o޼��"�E�s�X��� x	�b��P�Ҿ�S�^Q��m\�e�҃���-���T��wKw����>݈`�%���ׁ��v�.<nm@K�H����|�U��9�rC̵];<P��X{M�۰5�!]N)E Ʉ"�*�W�~'��	��\��'�4�j���x�F��B�Z$h��8:ҘŨ��I���ږ5��DiFǀA��Ta��Ji�7��Y��&����14���MawD؂	��刚��b�4c��*�\lx	�W�C��#1�8K�t�4�kQ̛0���*��ݸ.�hź����2���M�ڀ�'B�����Moτ&V�#\Դ|S�q�X/�}N�8�B�d�g��"ZS�"jT���ß�^�C/�7 y�@/}�G�6�!q=l+V\�z�\�?���z��j�����z��'7�Ŗ��w�����c����y��
����7o�nf�0�
�4��6X����
@q*lS%�B}�e���	�lp�H���;B܁����d�����d��#̦����_K�-{ ����<��ԯ�Q܃��"t��Au����2�<�n	0�ܜ�����X��2QwK�ॎ�M`zu3(W]�Iw�QB������Cuz��bxo/?�9�{�xC�OG=^�*��
��ÖC�n�q'N��7F�P>�Y�|H�tu�Q JN%���F�D�H�q-'=p�n�?�{�)l!Ät<RЕ����V��o��_J���ϙ6�{,h�9�2Z�ɨ�`ם/�G���<{%W�Б#}u���o���e���T�cg((��bQ�Yc-���<��z񝓻�ݚ��g�J�#�]yu^�̖����&��]]?�������� m$--ٔZSo�x�q:*�q�f�+��dԵ�× 9��Bn�V߰���y�����ޕ~U�|1
�J۠��}/xuq������{���XZǙ-mmm�U�KH�^�-jƬ�y��B,��7?��o&PY���\~W�
Tgɢ�8l9{a����(y%�duu��#��b�<d9�T��$�1`P�{Ub�v�1d�AYrp�����_�&�ڏ�<���$AgNO?Z�o���9衵8��BrD<�#9b���׼�Ij�o,mu��LB�%dxp��c�b��s@E��g dP|||,4���坃�g�� �0�;��"}�f�&bCKH��9=vWiˀx�ac���&�b�W</��`�CA�[l���b��Dj�*9D��5Z�r�m?��)(5[	޻L�2z2V3�ڃ<E�"j?�k1���#��ڨM!ccD�F�^p���^z-�ꏳȩ1mUf
q��h�aq�Usl�s�*�_f��ԘQ�Q�p����~���*MlE�=����/��4P�A��]�k2��ܛ�c�����6�l�H�ډNXآQ���C�>o�0`���#5F�4Z�;f�媠A�ƇhɃ%~s3C(���"�)$p�9�֚�s�g5�Ė�B��mKzH���ڔSM�R���y���ɰM�X��d��lq���5����`o186��6����HE<�]T���>��1����u�����t���GQ��ꊷƕ,�}\�hy{��Eu��dq���s`âՁ�������04���|k��r�k�W2�@_ˡW�"��d��oQ>�n�*$n��t�q8}����OFyQ����K��{c�'���ȋ
�^f!�D�:N�}x�>��ܻz��\g�@�@D�4�?]�g�=�%��������X�bIIV����w��)K�ů	гg�3��%��,%�+ϝ�6ў��7�[�AW�zT]���lC3����B��,ஹ^w�4Y\���g�9�����B�("j'��,/��*�=�?��_Ф<���d�����I������h�"��ghfc�q�1V���yVw�U�w���[�E �Y^s�c\C�Z'� *i !r�s��%=(�`�PId*P�^�� ��S����;�D�|�_C,��
(�4����"_�/p%�X�&�$VjP� ��&SA��!;�I)R��MC>��+˻/�B��e�54b?�,W�V9��l �Rzyq�3���.�u��Ѕ8�D���j��e-JS�}=?��)x?���ꚀIi]9������@�ˊӰ��S<�={�8,m��e�2�>����9KZ�'����^���B�D��e5~�(^St��>������/<�K8YdI ��]��$(�S	+�{��F������V��s6ռ�<������uY6�p�"�2~w$�ϏG{���k���P��|:����꿟����x�? ��Y�:�tg?
����dt�B;�����$�ߤDg�k�y��r4߸?f���n���a�'k���PKJ��0\Q{.�_��$� �����mj��el&�Ps���d��ş���?�A�?��V2b�k�]爺Y����x{K�&l9�k�w�rV+�Qۅg���w���h�����H`U`h	�
�,�J���N���}��F�[���Hv�\t�+gQIKor�RL@��Y�bE��`����wh����i�R�Z�����,�C������&x�@mۭ����� 38���l��[S(�Y�+�!Ăa	�ˡzy�hD��o��=︌�t4��4Ə�O��5�7��gs5�t~=Y-���!�>�
,V��MK�4((PT.����d6�}(���v����ͱ��]���(�w����҃t�(����Y��%^����Y{��1B"x�Û���Sl|V��x��)J��8�(Ok�K�3&Dx�,~w;�2�Tg�.v�XВ�Gs�@�Q�����`GXq�!�1jC�0�y�zҲ����B�>�0<`�P�r�S ���*8 �|�	���褌�@P�ҸQ��*�nf|��"k��Y��S�EC���!~�� '�;�͙짡:e�wB�jRS«Ļ�̔�I��1�Q=T@���a��i\���ǰ��OV�~���,h�U�,2a��QuUB�. z�4:��-q�k�f�%�,�!�(c-���C���d^�]]�����F\����j��rHU73�U��ph��NZ)648����#�3������#Ɉʄ�ε�W%���;e��<��
�y�̟�������J���%e��ib00 U��>}8+�z�<�� ���D�$:�,�Q	�e�%�a�����扎.D:�H���$�Ο��g����^�9ǻ�����x�゚���ّ%�W9Z�)@?�kt�uۏ��c�|���̂��5���ѕӠ��g3)e�Ew�e��c5 ш(i�k�񇃗�����2*&FY��u���r��
������Qy��"B˨Z*a%d?tA�0٢ҕWL�]�u��tR�e��mz,...Êj���v��*9�O�$@��צ���F���79��d���LʱX���ʃX���vd	zf��BjD�2�KRr�@UnD����l���$)����2?���}_c���
�~Qs��83Og�
�����#�3y\a��t�J$�� ���|�v�P�I1�k/�wRl�P(��� ̽`�z��lĽ���0���ԵM�.7=�.��b&�
Uy���c��:xśoW�f�7oޔ~��;�6#��I����h���@G�Vy��=<[ݱ�g+4��A?��}�Bs�e$ʫsN�ꖌc��ܜ��tѯ��c���9 V�Z��J�4�ʧPcPZ^^��模1>�zm�̔�;���;޻��x���tnCϖ��s3���5U�B8<�G22p>�J�����&��Ŏ�}	�g�4~|6B�o��)��sv��?�����L#z�7�{bJ�|m�-��y����`qTB���4�A�T���Q���E�Χl�Z*��Β��u��4`�����^t��~xS�a�_?���LR��'��(à#�!=��8|�qH
dyͽ�-���?��#�/�$�u!�n�\_��5F��u��(;��p�[�q�W�ZP��E%#lZU�|p�8K�,��e��B�h��|��Fш��mTt�^�؂:�o��vQ���'�L�-°��ꂚ�jΙ�毂-( ]�O�=������xQ�A��FMz���S��?�K_h/��?�X��ʷ��^������T?�����Y�q'���#t/�-V2���[����:�oz�둃n�u�sҋ?�,՜���bԽ���O�n���(�d�DܰV�I
�
��y�y$5:E�n�M��n�)c9�3���%t����#{����e�r^6HBPȘ�[��q� ��}_c� 6�%1q"�W��b���a��.���I�7�z���5FxM�H4��Km*�[K��F��`;|��S����� _yZFA{����"�[hM��-6��|�"=({B��f�)���0h�����V�Κ��p`AG��#t�W��a���x�}k���-"�i�H@��.C5�G����ű{���M?�DéP{C�W�Rsh�;ݲ*4�� ����9�pp���;�+�����`C�"&���ˊ��ǭ���Ʈ��h�H嵈%k�_��(̛/K���
snG�r���#�N��.������"ȧ����a��x [��ڽ����.�{�A�l�#�:r�F���z����/'Dx'''SUQ��p�F��ù�n���Y��Ʈ	��`
Ms�DԺvG��*�n�gD9��,@�S�Wu��lZ���~�4�$��#.e(�#����@�#�m̃�o���8�w�+�o�^�,Ԋ������JV��]�.}f
Jyq,�k19Θp���h�o6ߩ0~"�kě: �UÊ���{����<�A��hʇÏ&��SH!5�������El����:6;�|��W���_s���]ZJ�lbo�S$�;�:�$tں�lW�w'�M�)5�>�Ozg�#�])���e�t�aAQ�{�3���G+�]�j�P#��Y���롣����v����GTi-UhE�x9��#��"~U�	��k��o7��fy����K��$�7�ht#����U�y�׀S?�M��}�F�_ғ��Y�"�6p'_�ŷ5}3mMr���dٌ���5ө���K��mM�3ON�(�:ce͊�[��F�IĦ�k>�ey�_M����谰�ؑ�m��͚�A�8z�^�V̊���m�k�3Ѷ��r?'1)�W��D�@��~�>B���,�%�o���=6pv�T�2����b$�DA��k2���_���?JJ������ʂLf����O�񄬯u�\����������Y؂��kH277ϛ�݈�
�XL��AS~ؖ�N����K�?��G��K�fr��,�w鉔�4�!��`�幝%%R��"�R���q�ހ9x==�6eےoP��2~<2f�N"��6#��"n��
��ts�%��N���q-I�}MFm�Rt1���=�j�4���'n@T�vU��D�ï'�U��M����mE�I#�.ĥ�;1�g	g��5FfcN��� �ڙä�=������������A��1��$МYH�`�Q��XnĿw��v$`��~EBq�y��,����b��7Ԃߘ�(����R����
[�0q����M1����5� f��|�F+؁<��ʯ����mm:7V������-'��p��q��Wn}��I��a��V~!�����c�ņ�=d�iiE��ͤ�E����C�[,Fo��s�.'.��r&w����!�����X��6�.94 �'ќ%�����e��~����>jT$����%�\E� ��Ћh�a�?$n��g��\(�>�1j!$�F�?��^�y~�x���+;i��[x��LFV��K4`9o�]���zPk��<��i������&O �;X(�|	��z��tV�3����3��O����,..~\e�/z %h�Es��/5&Wu��&�e�鮒]��
�1�R��N�&=�\�R�����?ы�b-���x<7D�����@}*�����R}����J��ʼ�8�c,�j3��6e��u���`� 邾�[���z�&DI_G��G����(�:}�Nu$'M����$z��Ӄf@:�E�8��먟a�2�]s|�nA�R�G�>@��Ȭ���N�o_u1��w��0��T�5��
�`5Q{f�|U.�Ýŏ7ռ�����3�`&���R��܆�r<�r�?����C��X_�h<�'�)�mO��.�MB�����VzW�vd��U�Ucl���ȍyO�j�m�x5�����|�Kh���@����T��D4Ĵ�ƢQ�y���S��a�g�ξ���������^�e��R�:ۆZ?���,��ɩW�N�=�0
{�e[�ji�|L0ƬG�MC3|6��f�$���n�!��9�WKA���P�{��z-��e�ѓT&-�q�u	\��LFX��|�v�U ��K����hs[a'��GW���<ז�M�+Ȃ9��]j����{���Ix���MR�o�ysw��[S��Ы���:��7�Ԯ������(�z���z�2&M8��j��?�Rgpk��c�i#�o��A�;"��CRs�yj@G���0:�ת�4��T����]{Kގ�x�I��ȒH+j?����W���]j��
?�v��d XE����X���&�<-?��e<����O��(0�Y�W%C��I�x��h�`��S�*ǧY���@����P�V<L�i�ȱ�co�Zʯ�k�$^��.F���r]��ZCzB��e�V{Xqsc��g�/��X�	��P�*}K����ѸWgu��	E�r�E�GVJN����:'��P���g?�ĒM�.�e�ؓS��{�c��'�Ю�eb�R���$\X��� ߘ����ɋ���x��3�k��K��i.9��<a�p���j�����������p�E���j�x^s}��NqS��ͷ�M�3������B��P[�B�����p����m�57s�d�/a�������&0e b�=�A��:��m@�OrHcs������/-�5ڔX���N�Z�%��{===�po�J��{���&΄&\:���.7}��c�ꨒ�k��c޽�Zv�9x���ؘ�#F���wУ�E�u���$< L���������QE9�D�gh���Ĵa�T�A5�F;�gU#@M���![l6�>!L�wG��An��6�"��u���ՙ��#���D�p.7G-Xv��E��i�3�y��8\��`ä1���.��s9Ҝo��6JR��̉�h�M�A�D��⭘�f��l5L.����n���݂E~��a���]18��O�4D��=���+���ҽ�AG�|�ڇ�t��n���2faսS����%�}8�U���?Mv&�t�$5��C�tOq���<�6���k�ץaW%"�Vr.�&w��S<�y	��MN�7���F���S,l����yF�I	j]�gn 9��懘30c�	;��=*|��m	z��y��<k���ݮ�EU|��� �ѽ���9[��[#�1HK+&zPE5Ҝ%�f�Þ~��y/���E�ԟ�>�������:�X���a�h����O�s~��j�5Yr�Ӄ��:v2�8,$	?8�idY*����­��.���۰]�0u�m�^z<%n�8�T�~ť��.*d�L��4;�i�=ų�;wo"��>�e<�6¿`E��t:��|��gj�ɩBzV�[��*�ʘ�����/j>�"�V	�+���vRB����ïo�9-��@����c[�a��ֽ�#U�^p�mWNOi`ݤI�gi�c�5�ҏ����,��dvǘ)V�������&�d'��P�MM�J\���B�LCл�C��+_8���%/ٹ7)��O���!�C���Ѡ�ȣ������@2O�/D���QSe�B���-?���]��Aס6��).E�i�F�!k>�����J����,o�FI[�$�<	�Y�4�-��4KS���L�Z��FW�GIKﳎ`ܓ��n��6�n��}?>G�#X=8gTu�O���3���^4�o4 W�z�|qgyAAiA�7�o��Z��e�c
�.�[[l���
y��=�e��?�
U	�s���2�%���F���_���Φu`t�K���2��h��w�6
V���P��M�7�v��;59�%�'���YčL
ee�Uk�h
A��Qw�E<�9�T����i��0a|���y9�x �=7irSqя}���� �Q!7^��l�k�d9�dy|�Ěw�7_�� ��/��e[�YI���8��݋b��'��5��!�q�^�C���n��D��'6��$��Ս���?xd��T�f���3'Y\��[5r����&CFW,�zd�v�u�1�	�&���]�br9��5���ۗY�Nd���N�3���jf�\ښ}�[0f7zH<�7~,�sya���֋�y���i�EX�
�|��OF�rZ�2��@��b����Q��K���+�����4�l�~_�����l|��6�ʜ¢���*7ը�r9
/Cccc�ؒ���3��20��P!�T��h\XqsG�	�#:l�f۹�_�g�my�����aE�"����F淌�#9�潣2����㞶�6�jY��w��'��������/v�L�.��Ųj�����H�<��9%��I�.@F�����vi�	�|w7)�fI$��ӂp|�.�A����S�H�F4h�"�*a�lN3���=�K���^�F�&V�{���E��KT�̡����l�nr�N=r�S�bC%wB�{�u9ύ�4�7=H��96,?�ϥ���~�K1T�<~�:�~���~�|��{�BKu����%p5ԉjh�4���b̲���Y�K㰳�j����EB�Hɷ�(��bj���b��;�[,��
�B��e|��;d!��~�gJZnV�RQ��,�K�b��&9���j�os��Nf��t���R����r"����t�W�3��͂�
� &S�!O��z�F��Db�R�?���rLf�D
��ς��j�f~V9�'�t��b'�Q����\�:~2�������XI㽋Uqc��mcs�c2p����~���7��������{S�$\���������� ��$�a��ʖ���`C����"~�1^/�HK�#:�^)����z#�?ni���(�o.��S["��ZJ@1�;)?�F��ա���\�ڰN��z�W_DIA��bT0�v�d�R���O��%�B-��7�0�O�&�7:��7��ʑ�y^n���4U/��EI��v?��"�F����z�,�V�i���d�Һ2:��P����kp�~��	:&"@�e�===�������q ����1���ȸ��lO����:�.�}�^~�	��)��j͠��z��{<.�4��~{�K�EܱM�P��'���S]óg~�Q;�=juGM/N����"���$g�^x��-z�濼6>������y�7��ԛ]�ۇ6$�=k�&#��ע�١R����%ɬ������K��k{i�E��c��
�{�::fe���C�?D�ע��4KRYO�{��*�P�2IMb�/�V/����0����Y���.�]��������g�`�����u�����_1��<4�w����C�J��8���?�^��h֩��r��I��K�` �cO�*�(77���S�jJ��I�k̴##|5wy\)!�}�c�A��)i��JZw��}����߿��2P��Ü����Σ��S;v���ڪ�a&=0"�6[�Sj'������z򑤒�����>����Ry�;��J�h�`85	a���**8�a�e?X��Z%�5�B���|B�� bg`��r���i�u�5��aY��5�R��&h�Ra*קu��>Ү]&p�tdSy5V��?���'Z�YDf޿��j����-*j��M�\�dJ��y�'*�� F��R�I�����\-����=��B�z*w��W[��]�h�KD�u&�9f/��P��ܺY�9'�I~����{�� �� t�k^�ʲ�-w5Ӻ9R�iR�@��-�#���&����[�ZFq3b�����ڑh��0�/?�������7P���4�V���(�4
��r�����Ss1����9YY�%�퇞��������1SX��؛io����|9������H�M�~�r;��ِ��#[�$�����������T;�a!c�#N��7WV��Ȓ���1����@Y?g�:3\�C����3�����Y�Ҕݻ[z*�W�t#pQ�����1�T�C��9�v��p�~����>P���o;Λ�|���찻�J.B�����}C� 6�Y�{}��A����k�a�8:&�
6�RyS*��"G�����������јڻ_?|�ޑ�2��{`��e�%��a"��U��f�UP�<l9�śG�E���r�1�lM��Ի����A~�\b����,L��kD�,t;k��23+�m�4�踁hh ��h\2Z�g�%�5�@|$${]A�(8x�Dvѧ���s���#9&6�̙
�5�K��i�,WEC��[�Q���A�|��̦FE%���kG��ろ5��x�r$N��iҥC�5�vG �s�\q�Q�Ct�(��������f�ju�2l6��Y�l<WM$D~�l�v��#��C�\���\<��f�}I��+*l�V"$d6BB�sғ���L~bJ��b`�W������˸/P©D�{�w�yAG��Tĩ���	;�A�(U^R�3��W�> ���f!�=�n��j�':y�l�ӆP \�3�k�(����<i�`�> ��8��.Je�9�_�r,���ܩ��x>�$q��ߥTb�H�������5�V�ju��������-��[�d"y�$�W�I}�g���{w!�<.���=i��>YK+�R`���Z�o��ā���o=8#������ʄ��ƌD��~�M䉏u��Ö��}�ld�ZzM�,TY}��.��x���M�����ېus���/;���u
/�B4�fs�,_j`2w�F��r8h��H�D�˗���Fv^�
ᰴ79!�����]���ŕ�ce����T���Lw�(��J�@00�Gy� �hv̻wUUUC���� �~,�2N�����Yk`�J�����n��e��AW�ѫ�]�{�����O��e�J~�`�X5���H���*��s��uJڨ�,�ٙ�}/6<���)��6h0(�^��1���)����w�mR-b~����k��q��6@���P� �~�E�s���5������qC�C�{����2�s���;jBY�$d�@֑��Ԫ�B�#
ɲ����lqR�hn�~rL���u{&�1&��e��F����P

F��#+���3�]3����v��<2��$�)��ʑ�{r9,����b�J W�)T��7ގ���q�������G���	����/C,$k��!�Y#�����qr��L�ԉx�VA��+'�={g p���ߌ)�Σ/��%"�����3o���|덋#�	#����0�H�0��JK�k�hǎ�VBfI��;.!I�F��a ��/5��h�*�D�7g��I���L�/,�#k�$@#w5��93�#���#����EPhd|7zb����Fഴ�Χc#�{�$�|z޾5�
�.��p�T�5�T�A��޺�o��BW�fNVVO�iE�p��H��L�}]��85v&�n�Cp�X�¦��CQ�:z�A4���@���g����N�A�5�����M�����"b!�J;���G+}o��,���!�=W<h��)�C��{z���;�B�f�TPtax6�N���a��"����(B터�7�EekUAyBBB�]Ʉ�x�W����f�+�ԝ1ۦ��%��e����t�J�"�AP�g
V͙���h��CT��*�����3�O��� RSآ�^"����٨[��p��0��E�Z˲���E�b��^���*
t�I����C��[g¼L��W��3��¯4�������Yݪy�C�iw,�`j#�ݻDk�y$��v�u}"�
O���ճ��BĨ�ii����g��l^��g�7/j8�[�Ré�ew+���c��*���z��&�m��r{B�nҪ�B��&��G�W����#�NOM���'<���s�"~ۋX����k���	!F��q�\�D�eڻ�D��E���f ��:�S6�6p���ߥ���)v"U;�N"W��O����Z���(P�R�5��^��ճ�Vu��&8��ޥb��ޫ���?
t��f����MoL�M%�p
�
ٌ� ����ۡ�?�So���Epwk��~�l�t������3|���w�;���O�J�,
�r����Z�9խ^���f�a�'/��ŉH��&%��+1��-�ǏD̡r
J�OL����z�;��۾�{��[Θ]��p�~�Tz���Rn:eHC�+�ʇI�>Me�gh�wT�nW������6�t'��o� Ũ
BՑhk!E�-O#<�6��o�]�հ��[H)nU��^�bE��W�&�Cļf��Q��L�}m����є�������68AfQ"D�_k�,J��Z0^����Jk�4st^�ۈI��� {Q;.swt$[��0)I�@'�~@E�M������=ܐYP#���e!"e��n�j�=B�p+	��>1�>sllLu/���#�pɛb�S�[�[��x�_Ղ�Ո��{���XT���hT["�p�2��B��1]�jv^�M�!
��jp���ۉ���>��r�"�"^�'�=ә����,Tk��L�)/8�Gq��7n�t���!���)**&m��4���~�&���xR�����"�����G�������L�i�3��B�N�<�ؔÅ	Ĝ,0cʝ,Ɣ��50�G�:�o�����"μW狋��2)Y�g��­~!WhN�s�{��0dz�HXj"]ZZ�#�3B�q�,;FD��ޕ�Å[�]�I�鯣����ۣ�M��?[P�No�D�o�`������5�9�6��Я��{��u����׷�K��B. [��ʢ�{���������7�$�xܕ��-8�:ˮ���s]V���.&��+|����3����P��t�y���"l)��k+l��O091�/rO�|�jFG��_�Y�%�Gs%>y���a�Bڴ�B�?����z�	�&�U�^a��X���k���5����v���z��[ii��Rn��9��91c,�
'��Gu�0��5{|���J�uH,p	�B�{]�݇' R�~,����_���sm��[�q#�\K?��'�n
N�;.f����|��0����炙p�ɯW���,vf�C[��pfQ�����Hv3��[(�MS!�L��C��z�=M��PwZ^��?��k�D/���Y���1o�Z�'3��g���E<� ��ڐ���d�dffz�F��KQ����+��U�
���K_��]JX��l7N�G�8#�0��l��>�M0�+Z�H{]7���"� 4j0F�S<�Wv>���
�,@Km����^~8]/0�j]�d�m�V�l��wF;�Z�[s������3r�3�
�����*���-F-���e�Sa�}��a�K�ѥ\N	��D�4��h6[�ڑ�`�<U��q�CĎ��}�î�ny�$����~f�$a�@g�H�����Hn���7�/���E�{M���Z�E.9p�fr��"�/��y���pW��T�[ȵ&f[������ym����fW�'������,�L���u
�Ի����s9ղv͠Yr���(�r\���[�V.����5�&�����T�&�TQQ��
�!w��Uy:3�kx�@��4��X��3�������E�F[`k����F������ν]J(u#�*˪9�Bݚ���O����c�<����T���3nO�Np���p���7��b<��RK��#7��K7^xl�uj��%[��k4~�j-�?_�~�TC�-Eƫ7�9C�̭T�r��3k�R�:�?79��W�X<�D644t%K�,a��,;�3���^�����5�:�7����>퀾��u��l��\�U',�X���!X��Z(bDP�;����
�Nܠ�t��CX���v��6kz��MM��=Q\AhW�4�O�~�80I���ϝN��p��Κ�q�B1��;n��P�v��]'�vy{?�&���O*�n�Mni=<�ҹ�p�UP���p�7ӓb���ct����F�h4	�S�ؠB)���N?�B�+�u���T-�J�[$5�qǈ�����>����]j��dZ�Ie�f:2<���k�B\���Qk��Ҧ��d��-/��·���
h�U�?%(�w/e���C�	�L?S�E���wޟ+t2d�졠�\q~4�ٱ��"�e*p��pښaG�N�i�����@��S��j��PM	#ʆ�'͒���G�F��nH�Պ�q+�)�@h���'s�s_���;�G �oD����1gRk:�W�l�}���p�غ?�R<����3��k6�P��j8W��-:�����+�C�����,[=8��$�h�ؖ��p�ȸn�^,s[e5��g��֙�e�����q�||�(�� T[�_�E����;���&k���4U��Pn�?[5k�+M�U;^��l���{N�o8�g�`�CX��ѓ��N�}5!�	�5j ��X3NO<�c�9i��j��\�ņ�OɇP���7���ۈw�D�����>�����r�:P�I�6�mZ��鋦�q���%��#�y��J���}11�mD�: 5n�D��\�~sJ3Yr�`iP�εx���6�����:��K�&eI�+��ʭ�)�m���n�RӁ��>��z��y��~7�v�\q���<��s�U��%�_�j��qϠ�ۖ��6�[��T���cT�YZ�;⛠��7���y�J��sw0(&�^��J��/x��G����^"BJ���R��ڵ�q�˿W	�{� ����ʫ��>=�^e�튩v�g�Tkʿ��Ӥ�u^��1��pqo�M*���2 Z*kMd/<�'���k!��~�0��	��@T��������X��VL�5�H##vH:Q�����lF'T�*���̐��X+0'��p<��c����e��(��;�3��ԋￓ�%�_D�	"�,�W2���Y����q�2�ǅfɒ�x��j}�f擕������ZN��U���4�ȩVB�;�t���m�պ�mfA� �jJe�r�̨}A3�� �+Gآ���=���'	{�	�{��"˔��d�)�s��@4�EH�s�����q���7Z'"�)���,�d�|��0wx�-���J��"���ƕ2����=w�0R	w�wb8z�|*y���WRS����������;�9�<�wu�Az����^O·�'>��k:����9/�G^g���[�`n֫OF�U8���>�dJ8�B�2x*,h�B�ϸO��$��ʶ�t^���0��ˋ��Q^[�?<;�S;;uF;g����`B�sK 4G*��׫ɭ�Z*�����"J�%����5�"�4�d$���H�����MX����٦S��~\��|�iV�1���d +<�I���p��LQ�^�c�Ff��������x~3�׳SH�*"��y��m����s?C�lXg�6�{�_�?PK   ��X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   ��X��g)�
  �
  /   images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.png�
!��PNG

   IHDR   d   B   �s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  
kIDATx��\�k���߻��d�dK�jA4F�H\BK��N?p[���/�C�P(n�R�?Ч�ҧ��o�@����UR�QS0�cl�.�lY�W���jwgz~�=������������;s�~��9�s�LBD�O�<�D�B�0#�R)�L&E�\��j�*����$bϞ=b�޽?��o�YLNNv���#dvvV,..�l6{ƶ���,�;*��!L
�{t|�ɓ'o���v���#d߾}��ݻ �;��n��������W�92H��I�z��h7"G�Ç�����HR^V�h���e?Iȫt~���Gt�#�l� �aQ�>�����C��m6�����F?�jK�Eİ�~�O�^����/؏���m��\.W&���������!���bbb�P>�o�V�#D���������
gΜ333�T*}�:��'��h�u��3���=I���b��	D��X,b���v!�o�p��
>pR���={&8Б�G�8u����ܿ��D��d)�N���3�������;�������"GM[1�] ��1��$ #.;�|�����z����N�:ձ�G��+W�xvg�1�T�P�����uk꣏���?�޸q�#m�!Q�sB��	�2D�uP�7a����;�B���MY��۷E�!�<��!��aw^y�uw��!��:>�!�t���'�����ѥ�·��"�Dx��dv����y�cc��4.=�����vD�t(��[YY���L:$ ����d��w���&����(��P[4g~��='d���.ҹW��&�v >YU�&�رc"N����0��r�:�P��ᡡ��r�cI"J�&vtx=ச���?9��[u��r�DMOOSL� cy �H�S͝0
�F����ˁ�V'����>H�#�0Hm�I$(��. �	��ras j��J�!���_��x0�u%5�OJ�*"0!���h���������d�C'.-/c��*O�m�ȧN�C$�.��:�UҖlo���˷b��ϋ�J�a�	�H�(��!��m^�0����͂���P�\I��!0!��8#T��`��ُ�2�F@����יt��,����BH�������>̕4��k�@�jnb����ٞ�(��5���`�7
�)!L4�
��2�'�G���SL 0!<;	�Ӹ�L�I���	�t�2Sf�~eɝ�a��`uez󃖄@l��4��4! :�7��,��U�&�B����4��.B�d�I�m����u����*�ج�;o��@�����J��.�v@�=��>h��@+�v�����κ�iG�:.!~e��< ��?M�t��ۅB[��݃��&o��|>��:jbB]uBM����9��J��!rX�"š��;�{����G��6U144$����V1�׮]���T�g	Q��TWu���ctl__�$!��q�������c/^������!6�����t��9}	�"��t��gGVΓ�;$%����~R}������{cjjꗃ��� �7M�����oY��3�.�:nCԭ��N�w��Mˉ������$=��e�))�f�I��`��X�G��g"�W�.]�300�aGgY~����_Y��� ǹ��s���]�X^��xNrT�K��xK�V�U���1~�lB�y~�h��Ż���;`�k\7�Ћ�Pw���z;�M���8-T�JKH3R��dB�`9-Bt��mZiK�XH���u��#=he����K~�/�-�D�W./���4�W$;>�m�����x�r@R5�|n���!����!��U����9�V�??�mC�H��u��W��Z�F˄�$��i���v��V;�����*�<���cx��6&��sq���"F�P��':�`?��OB�#BxB 8��<[Ӳ!��� OL�#�-�	���dI�+�I��ȟ��6ꬲ�V+��2	Yu�/Gk���5�!�kE�C�:�WiYe�yΕ6��D6��m�0G����=�>��C(���5ǳ�Q	Q��F]U���!->Hû�ePG㍫?Y��5;��S	e��T櫵r��)�#B��$�S�����E+���)���-is��CTP�Z��~�����6|ޟI�*"	��B_��7)��ׯN�<�/����9�8j�!�mB�0��Fj�-L�Q��8z�lI!vw�w�f`qH����fg��ŭr�r�5 �~��Y1���������+u \k����u�a2!��N�:�\�{�m�N)�D<�X®�˗/�x���m%>�QZ*�ga"{�&�JHPpI

+�Lf�}�K����و ]!!rX�$���Q3ݽ���9����SHR�I��%�7Kk��d�jB�3!�&��u��&�p�~�\i��E;�ʌL��l�I������#5C��l�oT
��m\;�]�����׌j1M��BB,� �
��8n��{���!�n&��Hㄔ�ٯݲ7^v�Tn�qJJf��,�?	��{6M�]��u3NȾ�����<!j5���%���p�-�M��m�	+�z�R�,��	I���<dD ĉ���P�\+���:�nW���t	1�.�T�R9�n�B}	q���|������۵bص*�
���7K�X=v}��P	�?l��v�l��k0xO�n�����Wㆰ�v    IEND�B`�PK   ��X�р0G3 �	 /   images/cc0c8c86-b3f6-4855-b14e-2ffc61d63776.png��TT]�6N) ����ҍt)]��]C%���t��5tà �ݡ� =�C~}���[�����w=�<sΞg�}�뾮{oWS�ŽGvW^�:

A

N�] �����
R��B�Sli�:�V��(��=�]TB��,�/
*ʝ��((Z���so���W4��u{E�m��-
�_y\P~��y���ϧ�������#

z�������r9���ǩ���F1E��v�����?���Z4����f��㮣�$T�nj�lf����O�"o��[GKwS�7�N �7�O~��o�9�����n/�DGY�F��͒�������=7+!�2�D�ظ��qpxyy�{�;�Ysp	

rprsps�9�@�N�o؜@t*�O=/,A�n�.��N4�Ϧf��O�����ϟ��m���%'�_�:�q�;'�?z�ϥޘ��)$���Dn�Ru��^���ĸD8����j�v�4uwv�tvv�������O�9��~�T��FU�P�?3$vm\�	EE����ԝ%lw��d ��{�%�^�F�(zy/�^��ڔ�3���8Z��>�����Q6�7�'��
7��5g�����H����B\�NK�N*著���*���~����a`�Ɣߙ�����R� �'X	����
�<�ŉ��/ay�`*�l١3����YT|�����A7�� ������pFY_��<��Q�\$.*��!�����b��V���	�]�hwOM�E���9�o!�|�hX4�(��嗆ɠ������P�k�2^�e���P�|�S�h��ҥ}_�NTw�<;K٦�{l,��k ��]��''��H���{���<��J�_q�Wea+�O�����x�%�0�"��e����"mý\�����̯���yn"x���{DX���l;�c����af�z��mj�N�V�1[��K��̂N>�:X��G���1�Ż��ޠ ���_r�{(�����'�Q!jY}�4�Q���?\pZ�<Nv?>N@Ak�"���aA�[�l�3ݿ9(hN؃)�W��Q����X�(�D��U
� ,�MΌ.w⊰��؈��Ȣc��"��l1�L&1��=`�����K��� �&	5��@��%v1g��3���>���3_Ͼ[��h���R�d��h|�)lM|`f���KB��4L����/,e�8U��-�̖�K��Ӑ�W_@"+����{��pu��z��i|�<I.��i���͚����F���KB�#����ن���'s5V4(>�g��c�9�WH�x�P��B���v�j{X	/iW��_F[l���W�%	��a�����C������wC3�)�)^�k��kD�-�)$�'�.�_�/|�����Iq;݋��+3�0s({5\������Z�u5��@1�W.Ձ�p�D�^}���b��C"��>�b¯	��y���w�C^�(�Q+Et:�9H<B����p���;Jh)��\7ߣL���w!��7ە�PO{RE��hmZX�T`Σ���|x���b;p�].�_�m�>�`��"�.�~���ir����P�w�("ƶ&M�H�]\�XeGD�#&��+���Iť� �0�f�^����zǼX�,���I����.l���`��#]dڥ���$V`ُZ�V7S8R��ͽf���[Ěe>��/�P<��OR0�z�*����j�=c�e����kBп�$�j��t�uO5C;�q2K4UxA�<���i�i/�s��R�!��'6�m .>���qY?����a�������[�����?=9rE\}c��&����b·>�+�g7zZC47�kʋ����37�8%�ݓ�6��Ѷ�XRf5SVa=C�4y@�?9Y��{�?y��T><0��V)=�0���w�c��I����iw9��儑uH ���ò�C�뽜�����fqڞ/��R%��$Mk�e����7���d6t�D(U�L9��^��<õ��"��2m������6V&�<6�S`���cǖ�5�S�մz���Y"1�d~~��<3y>����l.��+��k�.��@�@�P{�l���*��]؏��oؕSFNV�Su��d�3����UM�-�+������?$�=���j-��g�T��xSʅ���SZ�n?��@+��YU$Zl�K��*�\�{�ʷo���P���1&c����g��� 7�`��3��Ϧ��V[���i���";~�Q8=���V�� I�z�e�A97u���%�c������pEX�Xz<��-��"�5�����N�y=��()�M�}I�i|��]"[�f�c��6����$��.���
7�ܺ��"X������Q�%��7(���w=�Q����P���˹���Nh�d�s����[�y���8S�F���������4����o>uU��l3mLnR��Xmoα�����v�K��3N�H��)�X����VNa&��
]�+�'o6�?�O���oŘ�?�W�J�K�<D}k�Wp&�V��]��f�>BF�W�^��7��ybX=���a����^��n���p
����+��uSK`)���69ԈS^�.lTF�l�2�����b�4�[�ȴ�����_[��&E�UO��f?�$�7�[I"�OV
�zH#�6h�����qD������9v�ˬe��
ӆc��D*��Y�����!��D$��bţ��H7WO	7��?.������DV���������L��6!�PB��@�M"^����Pq�WY�Pf]Y�o�~3|M4��� Zz'�p_ؖYʲ��%+�!����{5Lz�l�N5���p�\"���ѻ��^�+'�� K^;]�~�y��zO�Z\��Y�k^��mQ�y�Z[g�%��ϷS��:��>\����i��r����b\�[��u�ݖ擢&��:@�9_���ɑ<�|T��g�	#�^�!r">��%�RB���Vp����t��S������N���?^ȃ*%����I=��G��$��=j�<ȵ�(Îs�w��*���5y�(Y"�E�]4 �1u�B�k�`"&�� Վ~M5 _tm{���.��J8�6*��z-.�:p��[���Ǻ�?/:�%��QC=�Ql=O3�pkD����m��5G�ýs�����x�'(e6���قn�p�F�u�z];��OsRދ<��
�6�W.�̼7&��7�<#@�D=@���Ʒ�e�FE��h��H��V�u�ud*?�0pY���p7�-�.��۞�L+H�8�Z�/���dAR�����阑
�>��rfO��L���������_O�g+8��1�v�"w�����z��{��O���d?ۏ}����wM�����ځ� OD��!�-��}�FH���$r�Y��t��.%�3'2b��"�h�(wI���R�4���%��t?@,d%����=O6Ģx��7穌��vF����7��J{�}�iB���U�A�[;��䌖M���'��מ���g�[���]�Mp TC�]5��>�Eߴ̝���{�ej�v��-�;�[{��l�쇭gF�yf��Ҝ1�i�2�F�?ʱ�HS�-u�{[��|!�\:5^���t�*�m^tՕ!n�P�2h�ii��U����as�<�9=�g?��lW�ߎ�R�(�b�#;>u򃢬�g���-> ^/�.X�8�A�l�}�+��N���Z֞�X�Ϳ�eNN��r��Ϧ�6���o{�7�ݺς��tvą�D�)�5�wΞ<ѹ��n��S:E���CPp�mK�7�]gs���j5���]켗����R􄃞�����x����;�����!Y�u��
������K/"��F�E�v�}늺�_ȵq΅�:;�z1!��K#n��V�t�F�;hІ�����11�1���oǢ���W6�{p^�=�7��#�b�.[�OM�:�R�<�o�i�G�Wx�gV�?Zm��L?1��у���B��lA�B�X�&�]v��{y?%�/1Hq��:Wp�-��#�ĸ��4�NFYs��ȴ��2����!l�A[۶�����a�y�
_�3����6��g7jV%�����{�?�hWj$-�l_��ߠ��þ�l+���w�ˍKw��q��L�M<��x�m�]æ�W�U��:��Č�q�^��f�@f�1mf����˶2�`R�E8&��i��`T��pф��5�������uJS��t3�H�r�˃��%틓,xb��x�)#���?E��OU�[��d�َMgQ�/�똃���|���l���KD;���/!�C��~1?dp��8��]�s�^�9���3�6��d̉�t=��tS�L1�vZm��	#�[P0p m v�m�QzDZ�聹�bmb�����&��_-R�A!�7궂�[��f�Z��+O�t��W~`A>�'8Uk��9�x>.��Y��h�&ȁ%�(LbԦ.У =����7I঍�S6���͸oe��>�Kv� AS�D|��/�B-m]A�=t�t���䍈Ր�-�C�&�Gy���S:#�V���!�ŀ��eߴ�e@����~t�a���j�7<A,?wDj����1��b����ѯ�)G�P&[ *��}bu��Lr�7�ֵ��i�5���oNd̡|�d&�w�f(�gG-sp\d�AT��/��=(�T�}A���f�i�g*$or{����l�(�����A�Δz�]gT����iB���gc����w�ϫ��e�e,�B�n�E��a�NԴ��N%���o�ى<�����Y�>M���'5trŧY�X;�#�9\m����+��ʊ��%�8U����J��gPl��HX|�80�t5h�W���6M��ϡӽ���!���,�8�E���yul�םt=��0�%�惏�KKd.�ٱ)h-�>7ne�2�|l�����&���w�!��7*?o�s�R�6R(��h>Y�6�l�+WV�M�e�+�<گRE��D���Z����q��n�i�9�ܿ�#�����>5"4g}��ug�g/���8?�b\G���X�E��[H`���]�:�k ]/Zѷ:\އ��MЯ(e^����n�^�T63*����1�/6b�>b��]�����k�xÈز��������٧�s�d��]ߔ�~��N@�5�V��I�A��H��l۲�5��D'�{���*����!�G�[UZ��=0br$r4p�A�1���!4J������F��b���^	�s�1)9q�ijSCc�u3y+��8�����	�y8���i7�Y���Ē�"�v #�d�V�]����3&�;Ъ�h�#K(�d�`�Hk��6yz�{�;��P�s���	I�W'����m�X�<�z"��}_o���>sU1���c�v�f%7��:�#\��Ure40Ӂ�E�O��p�0���^�O8$���)�i��.��L�ysJ�*�\���k�V
���bCR[��=.�N�G\J��)�xlZ�9L4��܄5�f����%�mU!h\N��;-��T&�7��l�K.|t���*�<�rfr�h̶1�oc�T��瑽�r �~��V]	�9t��!�����$����nh��>`��,A�[)��YVRc��2��nt���3^�J���ݐX�����r�[�U��l-�
lm�J�}=�?�4M5�3a�<m���xxVǗ:���Wr|f!vW�x��KL�Ӭ�kҐUe���]��	��E��K#s-��B�R�nm�WM�@�֖jD��̀81��hEd�E�5��엟%�<�G��{�O	��wܹ��I��t�Vk�xh󺲱8D���wkYηFç�晅��g�g#HG�	��GEh�ދk�Ї���n��xޒg�zƓʱ��^B_��l�*�!�`��L� ��͸/8*6�JP�;�x������vFe+x�'���*�>�+Y�?��E˶�Ѹ+�/�i��YMfض�x}~�>�.n�_��[Y�;�k���$��*eL
c�uu>N�`b$���z.�p\��\}e`�^Q�#d��DJΙPJo۶̜��WzWN~�?}�0�լ�<�H@W��'(�����G�_E)����o��Kg���%:m��^�h{��+��oP���0Qu"�$u��� 	�V�h��j� ϴ������xĊ_���~s �K_�gy��	ɨ�qOr�i�FXA������6�"Q�o�ߧ͏��ğ�8��*|�Z�P���{�~����ڶ����g����zW}i�0%ۊ��:N�cj���ߦ����D����������f�%>��Z����>� �`���C6#`5��+�AUwn��w����]�Nt�f�8<Y��^�v��*2G���J�;�x��u��A�o�E������2�x��)���]�b���}5���~$m�$�f���x߱�٨H�`��&p�M+%�+�r)��Q����\�7�@Z�'U��&;R��s�K�{��c�����v1���F��[�2�T%�8_���|��NN�^���T
��ƕZ�~��Z���6/���rԁ��<L/�����PE��&4Vl���y�UL��1���&|�3e")���Y�}�M�1�E;D(e׃̩ �-z��in�ǣ��̸Ñ�I��Ƈt�8XY��8z�c�q���W�I�r�P���B9�+_o}��Hp�Q�@������x{���޵�[;o��:���yͧ]�}�_�l��m�PK1<�v�{��F� ��<B�h-�h���$5��@�@�ɇ��i�Ua�x5�!b��'�k��g61Ʉ�;�㛲K'�<�N�a�l=#ě����~q�v���p��]_��'�,��`�|����F�I"���~t`�����)�+^�VX���63�%"4ߜ3Q��۟M����{�m5H�v��M]��~��/89���hK0"l{3 {;ɷj��,�`w�A�s<��p�1�3>�j����:t6t�ğ`.���3��5JxU���e�+��|�1���#o���n��xO\X��!�`���B��5V�<:��y�+�n����l:�i�N3����0���P�O�u����~#��v��%�R!��j2����0Q���h}�e�>#]i3����GN���}���j�ηY�E[�|�qҬ߇қ�o ]�.C�Om���\���	�{�|L���̨�f�|UO���o6�FE¹!;�r+scd�y��+�	''%f@(哸�L��x+{V���9������cT��G��~�K�PC�yG�675q��֏W�c<�{�f,s:a!�.��\��C.��|�ٿ/��}���zŁ��ŧ�J����{C{���v���	��-���1��cX^�狫�}�M�|'�b&�^JzY�mSj�����p��Pv�l�����޿V,�M^�"W�B�g����*	�[�O�þ֞1"��4
W�S-d�Y��Ӛ���}by�����^ ΛP��y���b�|�� rQ~lFh�=���?Uy�܌{�ѓ���~1B�8���r'P�m��'�M���~>�?�M�'�E���2'� �2��@�i�O�m'F��,`���+��	�@�ͫ��(��ub�c��eX�5��>�����[�+|�2FM����
6Z95����|�vV!��$7�'�hP��	������+��T�Yv�kz8�xu�k�R�!lg1�^x�(ac@��J0udL�d����ϭĶ]d�S*����֩�^46�ߎ(qb��55� <��˔K�Ԇ��]��Q�K���V����z����-;��k�(=f <l�0�n���)A:aݑ9�_[�k�d������;�*�j\�%�O�f �;<�r�l?f�v�9���M )���AIC�A�g5G�]q�Z#B�9�
wՕ�TaXSm�ʯ�g�H�e�������4�:z r�>�:��L�ki4��h+�J��'|�����v"�����s/��BlUU؂�_�;�GS0��_��Դy{�9����(K˒�}j*(XG�[+��W-0����-��l|\V�V�w�\Z��1��N�S&�8���7E�ʧ�b~{B�[�3�w��Z�A�6�fR+SB:�����x?�<�Q6f�R����%wq)_ݫ�d9��d¢���~���K�O��5��q�/9O���HSڌ`m<�9��Pw'�����G1!��l�#Rz/�H����l�x��	����O�e���EsM���j���2���c}���n<IOph�`��9�4!�.k���n��Z|�j�]�%%#��+��O͜��1��x�>/��<]v,�i�Yq�QK�C�&I�J݄Z���E�a��Z~��^��>iN�����z	cĳ�9	mО��!_���O-{��T�O���m�+A���6��ƹ ��HF��H�QlB���7�=d��W���$�X'�򗚖ͷP�ѾW�b���KH��Y�).�)H�`v��s�����o�>�c�����K[�	=e&��3Ȓ�8_@Ė@~1��{Q�!9$�x�&z��R8�on�`��I�D���e�C3�a� #�� ���
p���\�hBµ�g�������{�Bu�K�>� ,QY@�?� ��!�M~,��G��q��VELh�'���EB94���(*s��P�p[ �����O�ͤ�O�?��C����iӖo�W!=[�z�\z�s�T��(�@�?���Pq�V?�_v�//�ʗ�*�ug���<$�jSm�6�wI�-T�dRZ�Q� &ϻ��6��yu�� �5�o�p���5y��o������B��;��c���w�Qw�;��',HP��-���|�<�oB�FQ�������\:�Ǥ'(�R���M����GY��ٔ�t��u^LJez��A�l8%6����ɫQ6!0�C�JD:��u�;U�(F
� Y!���DdY��Wl�.H2�0�n��>�.�׾��OlnjV��$�d@���P�^�VIE�M����6�h�	�x�%)��2;+�"���>�V�م5L�L^���Q�P����		b��5��fD(O+��o�[�4^�j�<3�k�|�8=�>�x/-q���ژښ4�G"\%��������������+�~y��;��~�R�PQk����1�ם�穪#�Y��0%˻�u �Hh��o��:yJ�甍m�&���wM{�!�����'�X��*SN��#^w�4�yn#\��V�.F���G� �+���$�w���+�EE���Dhtn�E��4�N\����_j{Y���ck#�ʕRE�K���p�Ȅ�m_���s�e]�w���B7ѝ?/��4��x��+S�:,�	?�XG���-2����J��-��2֝��f�h�f����S���ێ
/��x������3�	;2�t	�eћ�Ɂ��ڈ����������dc�co�Yf��o�A^��},_�[�_�,�6�9+q�6�#+ �#5��vB�/�̅$�l��D��SF���l5�l"mVw/	�,��U�f[Ч�;��<>	W�b�	��/f9�1��N�i�a�(�`i��##�5ů)�;�����M?�a�"��]*�\J��Z`9~�ށ?�m�������LK��7*Fp�9 �F��}�2��5B��͞�β������i6%��s��㷴ji�f!�(������n?dp�j�8mOT���Ç@&h�!����L2��M�~%Kzr�xdɀp�ȽpAe��̫5�̴�Xt0�6F��M�&�U�~pQu��b$f!&pcpc02p˧%�6�� q� �=P;`�It�����E������.7o���W'P��&�1|P������;��$��KW� �LGv
>���K���N�v^�a3�=�Vܴh��I�Mڷ��9�|��ƚ6��6d�׷da�s�e\>��(+˫!��xJ��+�5�&nq�܁e]�!v��}*ɨ��
Ùb"v$R&pA~�KFm�B!���8��j��K��������e:�5���8%~����f����[�tV&�B�ݶ�.b,�y{P;��6%�ȇ�g�9�c7��\����5�'9ox�U�^3՛��!�X��'/����]��Kunm5��t[%���#=������[˲�@�؝o�������� D�^�OL�ѝ�<]���i"��.���G�)�o�ό�S=�s�w:��ׯ����[���p�X�S����,m�b:�7�Ƒ�A���sF��-mz`�����+ �����s(�χ�"��u�w_������N��b�O���U'jKTp,t/X�4�7c6�r[9�7���%wRK�X= �4� j�-�Y�!s`7�f�KL�@��7~�Y<!Z*���m���a}��)o�cm��ka�9�I��<��b���[jI[%%�A$�Gr��W2s�˃;��rC�Z���.ܵ��CYWl*ԥ��O7)��A�r��w��_��2�����gjI���u6�3yYn�͂��z�FK[̗#�.X/�=��"�e��n0�.#j�>��S3�J=�$��@�����%�kY��ƍ&7C��kנ���(E�y_k��{��:5Zٶ����4%z�xEOe�y��U\��9w�1k�S�l@7��K$�qhB������%��1pa%�@J��#�����,�']pu�9�"��]Web�O���B�pW�qg���vi����Ş�I
��=��Ҩ�"p�y-�H�_��ԥ��K����ZI�^��ʪ���<��9�H,ڥV�~�!nd�QI�G����]�\}��m��9����NU��X	�h'~���2#e,�?īK$��5XH��oݳ��%�e�6�
CR�ݗ���'E������3}�aQ��4ɂ�nׅE�(\l���'R�뼩"J�M[7Q3Y}�$�N[`_h�U�c�zGԨ���ŜO� ՞6y�oȴ:o�:�Z>�7��GC������C�3G�pϳ<!��bO�Q���owg&YC�ע�I4��~4x����~�XW[�3��Q�I� �|��g��d���芩�ߏ�G�)ǎ��o�5�o��$��k2�'��ˊ$Wv�.a�3Y��e2�'�19��e��O�\��K�"_�����F��G�
�F��?-P*\���O0�XI��N��BIo�(I*5���@B���5b�n��e��߇�I���͜-��r4�%����f�A8I=����P" C/���T�e��֬��L�S	�D�'��m�'�����]��3�Z�MM%�<0�/�+_l�mO7�� �nU�I����O!�܎��ݪX��i�q +�����>���ө�V�|ʙ
>��q�Hj���Qse|��T
ՠ�P�b]g�lb)�cu�b�^''���)~#�Nn�=����ozR��a��%�q�e%���m����uF�`�Uap�?��$H���oӜ����Lx�4��K	)c��ޡxQ�q"��^�Uj��f����b�?��^�]� ��Y0���Ӟ����҄L��334N���-0o��Wٔ+�=X x�ӟ�ɷ�xe����%
_���mc6����d2Ӝ�G^~��w&���jPf�y�F�{��]�ktj���df�?���:����U�٢�᳘����K��-�}���-��n��Q�U���4�S�/�!x^ξzLH �*$#�0G�q	���P;b��D�<�V��|����xn���3�t[��j���:,�n��i�m�V��n�\]���'E�š>pK�~���n@:�d��T6XX*����6A�F� (���a�&S
���)�)v֝f�_��6���;7ߪ��8M���X@����;ɾC� {-��t�����jv.D%����>tSK?zZ�8��V?RX M���n���'g)5��>:�e�*��ǚ���'�!6�8/-�Z���)�%�J�	�BO~�3S]&���-,���6X��흘H��?ռ��.K�1C�Tz��X��
�~�U<Ե�J�]�� z6UU�eVmB3�؀>��u��u҆N��x�.=lNL��Hj;*+���I���f�֯�P��(���,Z?�7�0<Q�#�Z�(?>��WgU�Xh�Rp�$3h:��vN,���CZ�y55d�Z�!�Q�K���a�p�:��G.\[� ����'��^o��L�S}A��(�L�0�d�5�%t���vFn����}�t~� .��>U'��������G����_�l�������	��X�� h=5�_��NDЋr�[�p#]�,����y^�2ޭ��71�m~���6�sa�5�N��[��;�|�ȩ�4�����O�$��x1�*dp���Ko8�Ra89��~.�T�/hPS������[��s2i;��ت|7�"}p�k8$6�D��p��� s�H|U�E�#}�B���-%̲���w�~����R+.�v(��쬱Z@��e�e(	�V�pc#*װ*�B��YX�������R�X�UUk�%�͒�?D�C� ɥ�#��Е����p<g�yx/o���&[oFS���D�6]r���d�R�?��Y�M�W�1�ʖ3�Kf#���L1Q1Z��~4$v�%�t�r�"OwZ�6莰#I���8,���9�HO�X@�N�l�^�x*�"�j��RRP���f���34����TCÄ��㼪��#�8ߎԩ����Q��~H��U��+��F����P^���f�#r)=$J�CK��K2�=+N��"��2SD��Vu���;�	!=�bv@�s\�L&"�
�֭��Y�ek^ٿ�����N�s�NjL����i�S.��[��Fj3"<>x�'���LDeKʰ�k���#߲�ˉ+��}�* �ekHf��J�����T�o�Dn2��|S_���Z�L����I5K`m5���L�q�^��f6PIm{�o�UB�'7��Z�b*�cٶ�~+�Iu�����\���Θ�X~����a[�&Z��ߛ8hH�"{�T+P���.�4_�1k���Ie��q�n<҇�T��s�v��Z	K�?����1�7329p���rߣ)-�N>�3o�)�4g3=� _	O�#%��ң���i��np��м}�;׃#IF�C(�]�!�!)�8�ܜ�X����P�OS|�!� �ab�z�)�i��O�L������<B4�Q����F����r]�������kզZ9�)���W��$�:Z�Mh��<�,�ec��#U��	k����@,�⹧�I� �4ֆ[�2�V��uet8η�Ƞ�D�D<]'�eno��-*��m��Bm�p�8XN��nD�,�<J�rm�(�x��Hn���NG��E�}�]�!�|��_�ܞԉ`H<��T���'ʂ�x���~?��*݀�?mP��a��zkX��]L=j5�M1Jpyi!�����QNX�&�ր��{��j-����X���5���pg��nd^����Y�+�1��vN6�6�n����.���\j�E�]�?'��,�M��R��<�X;�����*?���� sɁ_��߁/�TP�����]���\���>�d7~�����ׯ;�����q/Z��|0*=��%��F$z�	�;-�W�ߺ̂�9�Z:��,��'�'���&KU�=eմ�Ɂw��M�`���;̦V�� ���bRI�^�{�K/��*_N,I;�Xx�~�6�
�����:�B�9���Ӝ�dGV�<޲�h����j����¬K�vM�ӡ. ���|�6xA��N;��\���8��M�ٱ��R��M<va�!#����bдEnk���� ���w�f����N[�Ȯ��!!����֘�	FZ�����?^�G���0V.��}| �ft��,����Nɚ�w�FJ-c�:5�q��b���z��}�ޠR�7Ç���,������a�a11l��f(AK�S���$N�{{���5��/?�8nͷ��?p���t;�ui5�Y����z�=\� ��ۀ^[ڟE��睽|f�[Oa�<V0�����O�F;��
(� �.6�
�=G ~r�<�`�\�B���}�俹�����{�X�h�^���L�{i�(��O�~h��r������?��O��e��ڼ�|#�x`az�p�9|Mam�lay�☑;���_����Bt؋�2�g�vou���~� �1k�V��-�we��!3ɔ��ܓ���U?zp�-��`ۼ�i���lS�r�k��*���h���������bK���v�,�+S���9��D0�����jŃHJH	����'�m�)V��òԨv^�P⁈��C����d*��Q�Wt٢�/_\<��⩣�͔�U �l�S��Q�ƅ������_Dc\�����k��˛�_kN{��*����B�X{�F{y.r����*/��D��㒾��Y�J�:��g���{Z���a�7z�`���5���]���O�{�l􆆜����GKA����.,��q��� ��s��j��J��r!� !>�Ⱦ��z��_VyI
ދ�)ߙ��x&֛4Z��߽w$�,�(�h9.�v{5��-��v�ۖW�ٵ8�~%W*�9"U� ���o��![�Er�vz��29,S�RF2��g���*S�̽C�=���!.����(l�Cm�zf� ��Ơ���O�[!y�$��9��v���H®�.�&67	H��*Jt��$���xXC ��!M��|ɗ�>��`e��6$��8K����e}4��&Ͷ�m�cD��D������S:��N,����BbI�`s�?/�ɔZԪh@�M���W�P��"��� �$���ts蟯��K�t��=�eq�h�[TJ���w�8�bL�CoL�1�ҏ&9$4�.36�0nl_�Ħ���=~��@�郔�v��{�[m���µ8�1����|����ؒ�s��w�+��[��l��5��B�����FC[�YD�<���$[��^u1o���/���wº8c�qڬ(�-��#�(y���	�z0\��z����>o-7Qւ�Ddt�8{O,���óT�l�q0b��\�^��6#��s� 3B��1�sI�ohRɚ��cMN�����D�R��~�T �p-�u!�#U8�c���8v���G�,�-�5�A���W��5@��݋SkZ�i#�)ghG�sb�U�v{�Uwd%|���iQ�7��6����6H�;$�'���6�O���S�[�O(�&����Т�,F)���<���4�7$��u���[���� ��_�'�p�-��N�;ի�hjT�$&!�e��"�y~zV�8�$E�A2ٙ�'5�V�f��������Z��VN�r-6m��UߝO]�!�8�#OH���q%�3�!}#c-O?�� [�#R/?�6ܠ������G��՛�3�|��Gj���ˌL�������F?H���ۺ���@���U�G�IE⍉�%�������ơ ^�D}a��s�w9�hd��Z�B�b�T��3i���>m�A����>�����!��w������5/Ҕfj����bڠ������槽��M��ٻK�F����e\ID�d��m�d��3d&g��W!ls�T(��ϳ�z�����#�TUm�^@�q�|v]�����$|}�7�t�@mEq�]�Ý;�Ǿ���Tc ��P�C&�[Zb���ȣ��d���G`������1ߊKH�7����G+�HC����#��[pj��
�yvB�m����#��Of�wȼ���dR%�Y���k�99i�3��+?.o��Ĳ5R�.��w�.��;���J���Ǿc�E��'�Ou�t��@�1;��?�@w�9P�������3��h-�+}G�OoYC42W��m%:|%m'e��]�����H���Vpl� \R����g�;��HQ�8h���#�E�f���(� �2�c��Qr��U��w�?��(��3���
{,�_�f��F�	&��w�~�3�F.7�k�&Pַ��QBs����h`��-H��X8߼yN5�oߢѥ��p����)����5�*����D	�-��w�s�F�wψ��̹���a��UM�l��t?��[�IC��
b l{��B�tlظ=��	��lY�,d�zpI����+�G�U`@h�p���Ib�= r	:I��=zZ��k�^����ϕp��"�A��֖�]V�Y�#��J�97���Ju櫷k�nտ��mKW��/�G��0��b[cs[?"�p���K������`=�M)�/Q����HB��*lc$��'ۉ[�\q$�������B�oy%���Y����}D;�G�@��Z�u�ԫ
�F5K�L\���4������񥚟*����|�a*���6(������w�Sꢄ���8y~��jl��ׇ��ء��[��{JԱK��2�2}?�<���L\	�I�����Y7%�L�FS*�)u �?�կ�1	��ge�Ab/��W�̫K��Z���i�Pf4�xr�I���|!p��"M�-��w�\�+{-� �m;���P����S@�K?7Ĥ��g�U�M��H0�~�ЏG������ŭ�*3� -=��/��?xSz٢�a��0�v>IՍ���l$�&*y��])� ApD4��N��5�sʌ���|�X��s����׈E{�er_ݡ9� �r�s�SVOY@'�xT���ଣ�>mpT�s��}(��
2����w���x����W��uM��V�
�S�Ʋe��5[΀��3�=���4�:�mɀx��sU����D���2��Z�4�]#I�_#�|^v���J=�9�h�{=;�k&���+	8h>To,TY�L��q���)2��-<0'��Z���4~sr�����/�'��Ӭ�^����t�^���.װz�B�*�FL�c�O6>*�^��鹨���ݪ�|������\�}r*ёk�=�"zHķ�;���+�K����V͖�q_U���I���������}j�1U<憪�������D�-�2��M��١/�NO��p��Au-]��a$���@pww\���n�� 6������.�s��[oN����E�Zm��c��^����ǣw�g���QV*���>F�+�0(��ˁ|�[bw�C֍�Դ�;+���sAu��"�F�*�o�U~V�~�W�����=�V^1���r��XG�_�.Wb�dJ�������!��C��[m�9�96��u֪�H�V�7���&��χ��G�Q� ��.9��J�tK�D�eGUT������뎦���t���K��������\'N'���i������RK�6�`�����T=�W�����5�sj�jЅ�"hK��B	�	tY0���~%~�3m%l(��������ɲ7��rn>���e�h���YX��jta7|1q��mx���>;�:CU������ηN�C��K@s�����ٿ�㧿k�2��m��a*ޗ¤�i�;�>Ӂ��\h�X�1ܩ��=�^����W톻�:��Z��}��	 �;j�^�r0���4l��9H�����ūm�Nį��8�=��8hK�"�l��S*9� ���L�tu���%I��Oe<�����|��s�7��m�I�:��Z��x�F���pG�0"��Jxݟw��I���6s8?�����9���@M�;�NxIsp���U���k�N.j������)�^gEyRe�}��F�m���s.�^&��e�����6��j���O��t���s�9S�f��Ѓ�~�<Wa�&٭q	�}�f��N�Cީ���(œ�Z�X��L�\��x��] �{�n�Kg���t�L�nszw�yg��ϬZ�._Bn8yAβ@"���i&��-(YZ�g��'��T�ջ���3�~E�ǖ�]�M��2W���M<��g�d���^j{��bbWi����`���OPIyBb0˾&�,�=�:��G�
n7 e� y[0�V.���4��.��<�G<yfڨ3�:�7]ڃ��P��ʗx��b�bYU�����r[-W1kHS�>��p���T��-6Ғ�NiRɀҶj�!�~��SU3
%�ȿ�$Y"
X��)D�أH��mt���[�%�f��x5+/�� ӄ0�j9�d�͗�b�D��q*�t���q/�^�,��xy���E�/מ���^���������,5TFNċn�q�f���B8}N!�>W�n��(;͇���ʫ~�$i[�S-�X��):(=����Ţ�rq����F����^h����G6����G(G-'��hF�@*�h������C��a _�N�}�}�`�#$��顦���X�����)�U[R�)U1>��go�����غ�P~nB�ޭ%���"�3.�M�c�k*��Ic�� Od����k��`)k�� �GzJZs�hے�N��Ls:~��7�PkM1\d��=���Д��}�m�%��Pc^D��;�3�mJ����ދ:��}����J�LHq�A���������Y�<�>�8����oL��6=j��6��Zx��#�
bm���$�N���P���yQQ��<�%��"K��{���{闍[��GɈ��KO�J�rq��[/�J�NR4XBy,�`�L��̏��,��n�Q`�F�gF	ZIRP��6�ku_6��+p�~s����t������|Bo���H���L~Dk�x	t^W|� �Ф�]��7.���&0ܧ��v���'��m�U,�̧o�L"�H��B�B��b�8m�&���Bq�o�F�|�0⩯��F�~c�@޶`����S��9��6�Y�_(�8}��ӽ�v��+hkA�����|�.��	!pVc�VO�
�����T�����%�8���Ij}i�q�o�������
�����o=F"4'�w�U��sX0���?�Q�*(�d��pi�\U�׀��<�wH��'�bw'���OMc�r9Њ&�������)̿eb��رL��qC�NFV�D��or�Z�O���ph'Y-�sVg���#	LTӹ�x_Y�n#V J��ږ�{���� W�0IU�����i1��w^�k����[*A��N�R�(i%�X�t+���e��z~�%'n�zxY�( ���TF��g$�y�^����̣:?-���7��ξ�|�X1���_�_�v���~�; �k���Ȯg��ɽ�A(��"�讦{A!L��hWP������u�������E�b-E ��m�2���˾@.�OK�|A�(6�Z�i{�����Y�4��7���S@p��@4C[�@�3sT_X�1"	�13���,u���-31Km��>��5;[@�jp��p�u�z�8k�hV��x�ϸ��9\����x�p:>��C`{���L��Mc�p遃�VXo�ݗ� ��uT����?V	�Ejc>��R09!��eWi�<�̙�m0+az{�;�����l�08�Z'�?"�����?�����@\9��N�~��} �s|	��].s��`?�5��H��&�N�'�7�UD%|��1[8ٟ��X���i%��g-K�L�G:u�T��Yq�9�~d�?�4��y��������3�u7&�M�5h!N������
g�N `	dL�Z9z_�3���!x\%L-&#a-���8>��տc�ř��&IAϼ�ub߃��dҎ>~I�?��n��u�{g�ݪ:���f=��l^a�%�����Sq�_�?u?�GE �Od��&vk^X��Qry�_\D��r\�r3�Y�*2@b���y�������=:�*h��bM[e�'ٴ�O�B�&8�9���|T[�Fjq�7�Udx�Ä.�D=F6NBy+¾w|pL��(���(*����^�͔��G�X�{|L �ch|�ަ�V8'����X3�̢��Sl�����y�����+�̎��a��Wۧ82���K������X�9�vV	0�(Ai���mU�~?8�[��2R��nߪ�m_�o�L�z�������pvp�Ʀ�$�����g�m�t�ੌ�w����- tTKb[[*�aj����	j��n��!�x?�+��q��e�o���u/�"'���1��XDe�x�;�Z�f\�L5ҍ�w�_g��ޓ��$|$����hB,��w���w���� Yd摱/O1r�!�w}�Io��*�Z-�=/����%�-��].ʇ8�$��S����oB���c�H�.��"��Y�%m?�B-`���ٛ���B\m��7��X�Ͽ;Ӷ\�8ߵ�`'}��"u%��M�ާg��	�[�'8�9��T��Y]ZD��f�æ�?�"T+��.[7n��̪;���l�qL��?7'�ol�US�'d.�T��Ƞ�7#�	r�yY쏖��/.aj1�!4���w��`�����/�-����k���e������̘�Fux�]�T�[�\�O����+L�;���q^��O�Ң��Q<��/�3���Ϫ<.��f��G�,z��]^+!���6��{�4����	��Ȼ`?p�3�,�O�|	�s�_��PR���S��- �b��{�`R�'ԙmd�$� ���yӅ ��zs��g��{K�ר�N�U�x<K�������ǔa�B�|/;�,����7��y��T�󦒶��ޔ����, p�Z�>{(zҡ�ˇd����q�O��5��K�������n8��{tW-����տH"�[���z����?�,��s\��zy�g��Y�+��J��dgRNjKagk�	ࣕu�b�<�Nx �ߡ�~�,��M�?����'���9"�s��m��ߠ#a�/(�4��w��s^$<����iF�HA�����L+���y O�8��0{tV��Ű�y���ol�v���� ˅e`r�o�$��i7��F3���0���T�d��W�Z_�h���Hr��(J~=S�[ -E���s6�M~q��.4>���ll,i���i�ܮ����8uqe�Ñ]�h�/��#_��Rc�a���VECS�]�������G+�M�i��6�R��93}���Z�ї'�;y���x(��`2�r��Ha�"H{h~��N#1q�nʶ��o>pi2p?�4.e�+Y��.B�#����:-.Nu𒲌������~F��}��S�L�6<�\�֒R��#����WR[�^$W�B/� ��f����ǽ��g�����n�ǉ멛'0���2�B�nZ:����z܋쓈�ض�;hq��P=�Η74P9 7x����#�q+�@>����&�Di����z���UW���k�!$��V=IO���~9����6@�����P�[Н}�l:��)���7+��V�t�����!|0w�HAu�%Cw5?�߸L$�-»(��=�V�K���G.6�ð��=XMV�
g�,�z\���ͽP;�7�8*OS��Q��4ò�4o���z�$��D��%�/�����޸k�N�Q����,�=�ܬ�՝��3ʙ�߇�&f2���<�:,�`_�����,HYōmm�'dW��6Ȓ�u���ˍ��f�\��AAK�1u�h.&|!W��TI��f��A)���mx�`ymU�E�W�?�{�ޟ"uu�G'��z�qt�T��!��8ٚ�՞��2���ߝ��u�5]n��Id	��rJ��k
���2L}�L:\�Dn�y!a2I�MK`�����[�2�A���|Ԩ���Q'ˁZF��z.s��ۤ|�W�u���?�ݕ��l�eQ��B	�%κ�q��VgR\�͓����YS5���d�뾅9m�S�UE��6�W_hmm� {�@�8^�S�O�~�$�����٥]"�I��%*Rկ	��+�@ц{�Ӂ�(�F.�o��3>K���>���qXWoO'BJm`�P����Qo�&V��^pqr�9�ѠM��*��(_���Xo��k[e�qI�~��֝}о�^z��� es���^�w9��kg�s��3=�'~z���?�K�;��O�$�D+pa���4���[�^z�iet�F����x��QI�`��
r��2�N��I�8-�%��;~����v�oh�θ��PhPl��B���FX�׺�����h&}���7�/gR��=�ٴ�~o�Ø��b�Ut W��nwK�7E�i$��u�'ŝJ<��%�R����k�w簓=�!� e9ԁr�����6��$r��6����"���zZ[�_ߝ��򘛘�`�;�K�d�H,)��fƔ���x���	�`�ͥ:�V��'�&�������&:��W��j2r��L��?���.���N2x4�����,PGmV��ivQ6f��66�����omU�g�Y�+�AT���g*v�:_��=�%~�NI��W4��� .�[´�TÚkޅe_�n��R�r�45p�_�}�nX�����[d�Ek�VS�S[��o�?��(�=�*$�K�a�\V�������wǤ:��=��52x���	bX�Cfr�H}�Lj�e���l�"Վ��	nV����Pc��J�*j]=龊���
�6�a�5� �ǅN�-�'��*s��AϖK 6�W���l���;�:]�!��/�!U�J[���x4'�iY[���w[�<f��]�'bx��_�RbkHU�,b������އQxy��z�͒���t?����k��l�Z�K����ݮA�?�=���Gqm�Oh��i׽k�*߹3����s�`s�UrVz�j��	������I`���(���u�A�z$����C���a�rR�f�u�7â�װfkr�1/hVe�����Z_��w*$��e
,�Wn�M����5��^�S�6~�$I,l����r\�y|�<6��lM*�XT��6�vC��';\hȳ�Y����hu��7I���$���	�x��"����KY�Ŗ3���_[-k2�vQO���� >�x��zBn��]U��xr��RկxF$NtD���~vՖ'd�J���XS��3[����T����0t����/�faA�G��γ��[�q�X/f�b��.��?��;�IG/F��6�sj��[BC}id����Y�R0]Ģư#m�HO5�_�8�.��;��(��님_�������������ů]�#p�5L��_��˪(�k�Y���QPt-.�:�]ES��[�ץ1ؘ�w����9f�#!�� ���P'�P�2[;��w@�5LΠw<����k�h�X/9��ٻy���l<N�?_ �}3C{���*;j�����>oo��ҍm%^��|�u҆3Cx2!&{�g�QO�͒�Hb���R�]�)G�P��=]���N!����W����	���T�b���8�ߎƳ���7u�w_��jऑ�wpN�1֯�O�=���(�����ť�p�5��Z��Y6�T�0�r�.���1M���{w>��g�~�_��v��'�1`��+���+I����$���9�������.��p��*it�����h���Jj����sWђ�D;p����b�k�����/ǭ��zN�ݱj�|Bl�[n�iS`������%�L��4��lm��KK�#E�݌�z�
pӛ��I�1�F$h͉Y?�h7#JխI��*\VҌ�;>���A��3����8Y����3�q���B
\�����)�S��V����x�%�蚲:p2J!ޯ��@�_&ؓN��٥�X����@����p6��+��K�ؖ���i�܆/�u�I2E�5������)ј��YV�XZW���Jg����FY������Ŕ'�b�kwlL�5;�ћڻ=n�x8黤D��E�x���f˧��ᴹ)�\��0ӝ��hWqFXԎ�q���R��?��4,���`�^��C�d����w�2 N��Y������A*lȻ�Vy{�f*�i�J�)��1��C2v��ᏵS�з���҈�o�HY��͆��b+)hг�--Jh�w�|�20$�s�
�N&�1N{�-Y�9�96,`n�M���r�#��E�$�K��xH��y��6��~e��WҢZ�ӂ�'���P��o�pZ��Z/� ӳCo�?`�RtECV.S����P��&G�
�6k��j�wN(�=��I\/�"�^�cv��j3��m�0-|`|!"B۳��}�� ��SS,�v(�]��)��I<RB�I��wD��8=�j@�Q��Y����Jg�"�J=h�?�(82�vf�n�t�1MA��q�Wl��y��!t4�\�v�����G�����b�OM��5��8����"�pS�!�� ���z]��8���BX6ӏ\s��7�Yr�<��V����<�?�@�F�b�:�}�W�!�Q9�<���Tl"�q6WҀyN����h3d�8�P����@
|�V���mՆʂ��y����g��t�}�{A�-O@>���5("��#Ьٍ9p�`��_74�U�����L�̀\&@���������S��W�����-�|eEt��6�Q���_Y�֜���s�߀�E��3�H%�c}����<A�áN��#E�M�ي����E�����7$�e�Б�r�8@��=%��柌Dvz�&��jn��Y�Lɲ���GU�pn�-<xW�o���ݸ�?�!�&�d����N�t������=�����`%�����K����S\�?�I��b�{�-�P�O?�>����"Œ\HD2���l�$L�A�J+W�g�c�q�HE�h���3O۟��BC�};j����)����4���&S�Y,p&p��+uufv�k�����#p+��UBqX��:lk��^��rO����6i���2�i��gE����i'"���9B��)�S8E�I ��e�C�v�w�I��t��H̭�\�S�0���ʯr���}3���@v8��F<l���m�/��V2�ąt{&�E�|���lOۄ�h^W߂u���Q�G�� �'wFo7 9�S,���åbt{�b�<�5��}A���/a��u;�X(��|;k�2o��<G�Uz��=�/��^���oP��`@�r8QIF�^��d�{6�������Q�{g������W�6n� }u���2���v=^?��W+��ns����VX�p���U�Q��v{���ۃ�+7զN�_�x/|��^\$�`(I�@�E+WXYJ�26��e�����HQ+�H���Uov:銧[�w��6��!��:4�E������Z&�� �;�ћ2R�j-Ǝ�Bl�a��Z��#�We�~G��~σ�@�I1��5���
·)�9-�y�vڣ�`j �k���XX���8#-,v�.�U���OI3���2γ��r\,���c�h[���3SS4��\#jр`�Ň؜��氃`��K 8�F
ND|�VI_}lX���G����9�����	�;�Y�`e�l������!+"��<���p�^ʻ�< 8
����g�v�Mc�P���} �g��?�����+:P����j�>sSU�lo�C�
�0��;d!�$~'=�z�NjE|O�Ѐ�g������xH�Ru��1��V}��9�ο�CMf.��8j�b��n��Ei��4r�����SW�?,���+��)k�}��m��&��b�G7�m��J��+�e_������}�s��0_¸�M
C�͆��a�N�r=zO������3OM���̱�M�i�����ֆ"���/h��!��Hs��B��sv���:z]��P�Λ�k� T����Jѿi�D==�������9/�
�����U�iE��H����gH��Y�E�%��V���>�ؒ�"���A��"{�ul�M/��&l�@�Ps��+&kq�n�[*
�D���ɒ�/feo� ��-��&�Uݔ�m7`�S*�e��iӆ���&ՠh���hg�47V$CCQ>/~F$�1
Z��G�aG�sc��`����YIji:�?�Z��ʲ�M�F�pL�~���/V���>��~I�H�?xN��[�gŖ7G���@I���� �X+k@�R8�e(m[X\| ~��R1�͐��!�ϊ�|v/Rnfh�
*H��x�N� �]ߢ��i+2�0�?��
�!�E�$��^���}�����T��@F��w����cV�E$!�;N<{i�L.D�fֹ~��)��dU�n}~C�'��������sr�(��s����ٝ�UR뤲�p�_ 9� ���e��QQQ�O 9}����|�����[��{	�e�=d����؁��I~��͐�����ox�PZU\\�f�2���+䆵���=��v�9�k� -j�HA�s�3z勒��E�^277���C���)�����ki�ai8t'��� ��{���^�	SD��+���/�d�*������7��@/���Ht���6��-�j�c�~V+2Q��Ou G�kl�T2	\�{	�Րo�����鹓vA��WR�[�~�-OP:|���v�q�j׫ko�o�������;��N���He
�����a��`W�}���*p����}������@E" ��2�n�=4E�0���M�3�Ǘژ�H���`�Ւ��Y�u��O�~C(�"�RuE)���}�)����q�k�:��<�~X�$!ESK]����=����a�G}L����c���
HL	���|r��K����r���]c��}U>��U���ﴐ��jTFJ�R�� [g�* ��+��|ƅ5��s��@�t��������bHX�R]�=���z+\�2������}��o]�����$J�Wz�ls�,�)�F�*��"��j�S�9�k��x_�3�I���(�3���<��Xk�wZ�*�0�:q�0�b
 ��s��;N"�%J�?~8�k" LW-C�����z ��Դ� �%�2��9�|P�q1��h]*9����h�z6�_(��QUy�3pH����jqb�ƺ 
�Rkb��]�z��H�vK�l��s?���{gb�`�������!`襌ʘK�╇�����c�!�����G���$,S9������K(��~v}��Q��w$2�.'�O�,Lr�E�_�����H��C�k�hֈ���7�+v#t�[��gP&�o�݅sɯ��.���SD��D��m�mș|����!��?�1�.�9�6���o��y���d�[��Q�~������j-k�GP�)35Fk�8���k�Ջ�ܜ/e�����|��;��� ވr��Y�7�R��,�ۀ���/Z������E�r>�;k��h��o�y��-)6�.����F>�"$�������>�yâ��m8D��E.�DJ/�n1@�)���2CȚ:����p��q~y���_|�p����sղ�OX����I���*�k��ع������9�Hc�տb�:�g/��SE��7�a�|c<��vL�����T�_�xR�����/S~�f&@ �� xG�KQ�@�-#,w��{�%�b���>�!�3�M��Լ��I���U#�ļ����+���kRA޼����{G��/�S�Q��+6h�.��J��|��N;�!��݀����~���	�Y�\`=E_Lg�v+;��nI]�������ꜳ����t���$/�W\R�PY{	�C�R���l�V������
�m�ƇF�9����v}>)skG�p�YeI�$0�  F�>/Z�1J�׻�@3R$����:��6S+�U/|�!�tP�����ޙ;�ϲ���YVrb��5��ؖ1G�RQ��Bۢ�&���d��,�q��5�T#f�p�;go������)��9���ooVaX4�*A�wZ�?��D˺��4�2(=F�>��Nݯe����Y�Ʌ�|!qi�n�X��E��s��G�u�����K-���Ҽ�@jX���?{k��!�����a�	P�Ö<����(g|U���򪌄a�F���ͻ2�D������k)4=�go�V����Z�m�?�_��y�.(A�'�`�)Z�Ml}oÝ���!⿭rB>g�0jY�BJ��+���.��A��}6���Y�%��ᝰ[ʽ(�6u3����*��JQp���o�W�7�ӑy	�!l���$�æ��Pp�e��q�:��R��4\�U��y�ܜoU*�+'�Yw�a`�Ľ���>)���������?R���D[,` l���Wu����s�CX7��'�\���A��ϔ	�54��Y4�{7z�T`/w9h��E�￡�@�v��C=� �O�5Q�!�Re�i:e����q�Q.b� U�gȞǫä���D|jO�����8&�i���E(�a��*�n��:)�r�����4 teeX��G��}��Nb0���nꄖ�����n�F���
�����H��������K�_A�� �.���}o�D�Ż��W��g ��w��
x�x�]�|_i@}������w�?#�Y|��6W�uN
��6�=�o�h�2��+ۥ�S�p:�KP���{���"�VO4WҒ�(V�
nu���H��<P�6����*��N�9F2w!e��0�j���.Ru�+W�kem�Y�]�8�e`�I@5E������;&�R�vY���\��	�!�Q������2��g�L࠮=�������T�H�@��y��&VwK��"�/"����4�L>.꿇Q-��<��c����k���-�E6Q���b}hn���Z�K��L$�7a�}GEK|����������0f
Ʀ�zu�������#>�j�c�&(�XD �̓S��Q]A�r�w��zo_$XcM��_�!Bo_�N^�de��E���F���h+�_������iAR	Fv��6U+�S���}#�fJC�����G�>��Qo��+:��5�Q��Ԫ�t��`֔�
�}�\uO]�a�&n��B�i\�;��O��l���H���m��ʵ;6�N˟>|U�e����d��J��I�B%�QR(�+UWK!]��p��E�G�@|���������6:B>N>���2`A0����l"RǦfA">C�&=';'���ɣ���hV�����ܼ�>�;m�K�̝�-;=��2�Oni��T�F�/�r��9�z�{�wS0?�����؃-�+�.y������~�̐f`f^1��j�9��l|�HHL��2�7L�g%�A�V��@����
����1�5�;eci_�.>x��Iv�6��a�����g?��N̯{r�e۸	|q0t3��ۻ�-~�B:߬���[ݫ���b\-UjS�S�H�cG4|*�T��qWov�����+��!��2f�㕕
�5:�zs��L�C�∹=���m޿�'�%p�q�}��`�f�泥����/������2=
$�t��/�?|��p�ϻ\@�_�.�;�\;M��I	�:]x�mT����K�̳/,��*���EY��!�[_��z�����ƛ��F�Bp�k�ߪRo�c�0~����Y��x�nMMo�n��P(��f��q�6������-�k�i?��/&v=N?��Z��q~��l�;�pRύ����WIHD���pi�:g��U�}��Z�K݉��26�yj�4�= k����8g*P��J:H��`�q�EƢG����&����/z�� �_&\��h(G0��NS����m�W��I��1>ͳ��.)-!%�77�I씾f�,ZQ��<Ku�\���![x�7A?�.��^�hU�����������n��Pg�)^���(���u�˥�@�O�Je(�zܭ��2���^��O��dy����\�l�`F���LP��p7IǶwO��}��P~y`s6��;���c��IǺ��S�ǆB��f\ג�Tt������u�DJ�*�$�l�r3v��9,*�sȞhk��z+���������� N�R��ͱá����AU�gM����WUz:L�@�@�n�2��	f=�8�*rԄ����P����\�γU�^^M���F��G�-����m�(@��!/�mdJn��d2'�~N<��muFMo����#�:��*���@
���	�f_q�~X�����3ե�@�r.,"��H����k�ĺ15vX��"������D���"�RO!�k3G�g;��e�AO�Zcks�ӮLŠ�{ש�N��[���������.bZJ��ɚ�V����Ld�w�{{��Q^X�ч"���x�tGM���^���pYa�ͷ�ޜ��)Ŗ���G�	�X[k�錎�E��΅��~}��06���z
�y̎ɓ�~��ch"���<N�HP~��/Y�c�R`�����H/ūI�l�{|�fڌy�c�@�������Ф&��.�n
�N�z����p�w7
�)���_��>�񉻤����z�)�6�f�"�`֢��B/� `hi��3{�ϩT�o�r���AM3C/�t�2������fJ�ť�
��k�:+�O��89c��^���]w��ci)��L�2:�XC	��w<��ܚ�j�T���O�E�9���QVa�.�rh����*\�]'�y�=�VQ�-t�`�T��|񰕸c!�e�(G�p�7�0&B��BL��^l���aLR��ӹA_�h`16ԓݖW�/R���ɧ�}���I�hq=Է?��j��H���.��w��D��$��?����.�(�ptu�vDAxi��蘢��p�\���!P$�n�I��@19�BF�	C};vNP���*x��qι1�D��?�/��V�~��o7ڍ�0�AI1�'s|����ށ�E)̯C��(8;�7���v`����X��鄌�b�N���1�{�:	�P*j�O��e����0	��-�B��d�:����8O�����z�KT|�P���F�Alv���z��1n|Z�+EWaiŧBe\���� :��^�nzS%��:�(�SIS�L��N��W��D�`M��}�0�Ťf�ߍX��8m,�8(��~z����+�9 (��b�h.��e��9WTI�������u���R��;����,S	j�fR�p�q����ɛ���[��nXbxN���Er[��;;ܘ���6���0,�󼥌�b@}$��\G���Z�Lӓ{�	���[~�;�+1�P���եIV~/S ��!O���^5�Uop>g�0ބ��E�q_0����U��`IF��╀��R�3	�M�a�/��Ѣx�Jzy��8C�B]{Z�g7En��<`H0`HuQ״�2�UC~��#��u�;�:�QO�����V�]Y�IH*R��B�`q�g'?����o�9M�Q���8/s�u�,�s:I��U�l_� �/Z��h|�L���A�s�&&��Ȟ��kOſ��T�h%�m Ǌ�E��-<Z
�A�H�����n�{{J�]��5��c9aL�;��\ k�ͲP�_Њ����gCQ��U��s���T�_�&�`�A�b �k�ܪjG.�G�4�f�L�ր�x� w�Q����f]�b������m�oGʎr��\�F��^�a��[e!��j)��:�&���c!!Ҙ\Qu���v_�wp����Q�uD�C���w�c_�i#�4G��Y�Gj3�G��z�z��KN��T� 
z@�|(�L��#��u�&!��ҽ�Hm(�#����Kk�ƽ�9�SQ�D/�D%��N��r3`��.V�'�oN���wk߾6�skn�x�5��� �n�˘?�>"�I,����#[q䡹��n�a�<%S����85���V�+
kCX���������g���j���G�5FS���s�E�d�S�kB��jJLJ���>�^��`:���TL�S8{s�5�[t���|vϕ��z�V*b�:��P_��,���:c6 ~KJ⦤�F��}���҅�Iu�`f ����E���6�z���R5D�G?�fw�ف���n*��U��ܱtV:�Hm*�Q}�ʑE�����"x ��IYj����$�C�p���O�*���Cޯ8?����F=�Raa���`�����Ȫ�]�9���*<�.�}ť1`�.^֣��:p~H�{�j��V�f��i�Ȱ�T	�^I��d��Wn�\MB�:�����m  ����;�'��W����]�k�զ�j
��/�C669Er~)m��ƅ�Blѥ퐆\'u�<��)��yZ�p��F�X���!��B�m�:\�>��ѹm>�ʸ���ޚ��` �ԉ1@ Y�l�j`�̳�v��D�R+�{��Vp�Ӡ��ؽ�w}7fz [��aq�静���g����`���`b�����J��򸴱�������Jn%�w�-	%�l?B�_��n+�qwo�S���¡n�R����bXt'��!�Y�o��}]V�[ �%H�9vR��b�PSc��l!4�a��.�M��đS�s��Eː���p>)�k���9Հh9@�K�ꐸ\�D��@�TǰH�?�,};xb3W����- �5�}�l���R-)ߴ	�~�|H=!\ʚy%|����Qm�4�����C��q�L������.�n�����y:�g��L�?�K����GH�]��W�ޝ N�S��=�l]̏unn%�	�$�Yaۨ��\L ���E�_�6���2�h3���؈�<�v_�x;LA���Pr�,�饿�$iY�MBBJ�z7�|'Oc:/ 'ZJ����
��ȶ�����Hw���3a���"��wc��.��tf��� �j���2��F���!��N��U���y, |�6+��+��d4^�]fԛ����Q$=�硖**�a_��=4欂�� Y<�U}��N�B�Xo����b��P�?~�G3݉�X:W��A�X�ʅ���~��9���_����w�aL8����uC�[_x��ȢG[wOw&���L�t\�X��pW`��9BO�=C(�ӾVvsO�I+��������P]���5W�9o�ݧ�����j76�<Mx�mPC����[�`���mqhy�8N��v���ׅc.w�w�pbħԞ�o*�:LV� 5@��}����b�����]�F)�w�r��W�J\W��l�����>Q�-�Xt�����iu}%�%�x�il��q���ҷ_P�C0�x7�zH�LJ��Q���I���)�J�]�m��#
z�b���
�t�u�?��!���SO��<��ȵTwY�vp��US�w��9x4�����������9�K�R��زCt�M���� #���Xq�����������
����F��j/�fI�s9���)'�@�@|��'1X������i?��7c��u|�Qb?ђ$i���UP]ҏ�Sg&�@`�s!,��ԥa�<��ٌ6�+B�[�e(o�o�
��f��E8�z���1�嚪�K��D���.�Xtt����ĥwOo?MFS�{�~ZzS˔c���vṟ�)�;�,�;��Ͱa����z�M�b��r��K4P���8���E�ɳ1��1�o�}еD���Р*=ھj��݊v�{_���\��;���BO���g�}@�3�3�xX'!D�|�+h�I�ׇ~`Y�R"O�/L��ı.N�*����|�!h���9OeF}-&�tf���Ntv,��i�o�����cx����|=�!F���2��K�]�^��eB�/��=�_���k�-��>�3p�9�}�;�c
�ku�4I(�����c�0 �q�ȭ����L��C!�畻:�oW�0ec�6ڇ�T�����/r�Ls�=�HbS��4�Rr��5��0�H����]+n�D��Y��I�F,�[E�^Y�u>�����[8�������*-	Z�X����ol�.@�: a�X���r�!&k]� �6�-B���`I�C#v�i��w�9�c0��[� �*�JK�u�V���cĤ��I���������!_ؐu��wd����CG�!�j���G�f|p�@�����2�_�C��b㦜�$%���6i2ڐ�g?�r�|�e��1�A\=�rm���up_�A|	F���?kY�IY�go粴�L��!8��4� �	w� !��܂kpww���>��3���s����|�Y<�Ǭ龻��꺪��[���K�5x]���p#��O2�}�}��2�(\%m�*#��s�V���!׫_����d�|��	�ocs����ܜ	�
�1.�2ԄoҐ�c�
��$&U�f�E�q*ϫ{6�3/����鑱���-�D�_�����BC%\Tj`�����
~�MM+�3�eg�vb��pކI��ā�*}m_U�%o='C��X>I����Ys�J-x�"����[��&��u�?%W��g��[��aU�� �Ф:l�,�Y:Da�B�=Jb��9������f���4��t$��ܿ�t ���[5I��?y��NZ?{y9%�^���զ����l$�E������Rr�����}�R���9����a���F��C�-GH�m�"֢x�؀G))Z=W869�f�ڼZ����U]����"��)��p�6���8�e߻E�*�u!\@��I1<O��!��z�{��{����ۂ�6nIWM��bl8�}IQ�8,�)2�O,ֈ��&�s��P��Ɗp��ײ��v��h�$(Â�lm���B��J�w>�4���t��E�`� ���G��3,ȟ4�����UK�!�z�H'�#�&^$/��`-\/����a�U���Q_9%����?l���/���4��1+*z�X�v�>��K�;x����ǭ�#�p5Ot���o|+��D�.�������ғ�Yݯ�j������Y	��ʵ���к���i��î����=+o�k4���};*%C�%h�t"J�0ؿ�NIZ@/��BƲ�F���,6X-D�{�OuD�����~{R'q���S��o���9J�㢩�w��*}P��쎅I�liI~D�Ig2WY����X����zW�hwl�!�+zޯ�=%�oCV�_<�����vH`��疬I]��}#B�ܺ
x���T���h��cZz��0�v�K�S`�T�_d8$�a�|�W�E{�|�?D&�������y��X�������)�d1)��|Y=.��(a 2�3�nkA�d.H�a� �wT��^�Xz�������u�FO*"M�SmӝY��mdX�b�v�C�ªq��V��s�o/�t��FHxOF�R���]\�x���v�|�Uy���~g���9�L����z�8��N�N-�Z�:V�ة݀�f�"L�+ނU=�8����_H]Lմ�̊+�nE{�Ed�)���CE)QEG��y�-q��vH�h�V8��Ɔ"~����fG���U�l�1��{Um�z�9��L���F���-ʹ}�v�c��.����7 />nn����Ԇ?�sy���8F��<��7�;XB��8� ���9k�/*�]-���3�(r*=�"��o���Ϟ��y�L������h.S\�4��������%e�����K��V�D9��ВPPS��~�֫Z�ԛ�k�u+߁Mc�����*��e���5��GBHr9+kh<���u�\�f���$K��[Nmg�l��v��o�ԓ�Z����tRD�)S�*��o@�d1߇8/����]�j�bA��0/��a�;,��|fm3qB�����+4T�"�#��ϕ��ii�-I���HEOѹcCX^a�q�}��s��!aTvo���ޏ���:4&��T���m��p�S �,GM�TJ���K��ahh�l[��~���"�@��?A��4_!Qa�����K)S��X�ܥo	���D5)p��8���n�+ƀ��*d@�����j����o�O �Щ��Hb�w���Ӆ3��%5f��ᜀ����{!F�n���[hg4cfr���#���7���-撷b�馜��;<]7j<�+�m�W�.k�����e���p_�������:�>���CKsK1?۱�܇!=a|q"�A�v�,�eh���b�
�����������J��@j�#�/�E"���D��G���U�'���ݱ'ՋI�]%KB"��>f<ս'<�l_��x3Y�Of�JPNj'�
�A��!51���5�[�M�n�>��d�а��썯�M�L�p�^�$�&��(%oӇ�����2�-����9k\��s���*���<�P� �� ��R}����eH]�,~�3!^$v��E�~lG�fuC��fT�Yj�2Yl�&Z��Z�M�~|���Q�*��뼘�QY��ṱK��
3$�[a���%-Yo6$m�'�w��4k�?���m6��N�S��1�T<>I��R}ǧ�rf�(�8��g�j��rK�a�|$XJ�t1���*�MH��C���<�n�l�&ybn��=U�\�N�y��-���DS+:ˊ|�e'��9�n�۲Uǽ�K����Y|<GZ��U�{��b���N��6�<�#ù'��R��ZW�Eu%�֒�p3;0����~RM��D��p����&�)�4c��N�u�t�1i�a����\��В�8�H�E����.���tXR�b�O+�k� uwZ
V��)1݇��� ��ןi�q�	����L2��N�^��A����J1(ޱ�e7�zQ��>Hs�{�;.�+I���bYU�����|a.1�smj�d��2W�1T�"`S��)� �X�ݶRoޑJ��$�~2wi_jo�d�����I�K���5��Ң�^D&M�|���QfcK�!g·[K��_/�8p�<|3��q�sD2�.�H������f9J��5+ϩ�)m	��m�����&�v6�
s5��V/�0S�p ��)K׸�Hr�2�lK�L��rs��L�Gn��܄�d	�|l�$�#��6t�~lr|�w(�J�cvz��i��%��tk!�8YS6,��2�Rro��+�cFK�A(���ہ�=��b��u��1jo����*�n1 �1�wy�A�>��̽_��f�KT��l������I��3�u��.ڃ���'Im9�@��s?]�W�翹 \�z�p�mo���N��9��'��R��/�J��
�F\����5�v�f��ː>ɧ4�$D�-�������ze�@N���i�����-̽Ey׵1K��՛�}̷��At,���`�
"rڕ�]cs������G�,��,��k��1��@�}Y���lj�����{Yc�y@I�=�J�̱�'�~�g	i��7�Әt�S�}YL[T�Gg��h %�x�d�aO�Ž�]�s��{��=s燺�hGj���%����z~u�!t�O�D��+ّE0��~�����S����Q��s�I̥k�-�5�ӒhMfG<] X�$��W�����z�G���T���Pm3W��݉�i=q,�s����R��Gg�Zj�2S)2���4S8�J�b���:�C�|/�>��� �l��/��F�x�'*�I�PX~�"�^��J����HJʍe��F瘂���ρg�+�ģ�/0n�}�ֽQIu�l�	�3x�>���I�+^����U)~=w���0<���@X>��Ӥ��؞���$����6�j�{��Dt����YԒP��Y3*x>|B�{}��d�wȥ��L�iX\�6���͝�m���^�|%}���^yP��$m��V�&����j�'����t��ͯ�[+����l!�=�&���Uܼ��
Ĕ�PV��a�m��aMni��D�#pr��)X�fQ ��X�\��I�0G�Fym��+0�,$�I'�ӂ�l�8{�RP�{���g��a~	sH"F:8�]��;�x�2E�|{�B�m�D!8~ �w���-V�h�lt��]�h��N���8�ݏ�D��T����C�Lf���)Z
ƣ�a��K9s�$Ϣ�+O���(&H�DWa��Ś�@���m�2?�f�z�P�Y���vk#yގ2pl�g6I����Km�`�?�<{/R>�P� ��G��kF�ٝ�@���o�-�+m�o[�>��������RIn����5�)�R��HEs�/N�7�;�<A��`��9���O �)"r�=���XJ"g �b� ��Ц�i���<a�uxs�U��Or/�d v"f�yN0��T���᧚���Ք�5�s�i�S�`�p8����+�:A�Z.�S�^Aj\Rvo5�*f�����d[z�Mʿ|4%h��k�`�Fh�$Q�N��כ���͵g�`�33�����7f���S�)��O5RZ>)<%��|�@8bFOZ\��k{ڒ�����4<z����Z}���J�`��xw���"��8�y5�=��o9�>ĺW�{]�d�\��V�>����ƴ�z9�b�v�D��n��<r��nSn}+xG멎�������'���ꋺ��Ҟ3����x0E��]��n��[�r���	���im!�;_" �FJ�3�]��}P��l�WÈ������:�0����o�6���e�O|���t ��w��V�T�N�.�N�Y��h�r٥�Mb�A|v?��|׮��	��/�Lm���i��-�8��>�����ޗ�U��,���HK�)��tΪqe���$��v?��̳�E�u]�ٔ廜(:���(��:�nHtgs,\�0��'���
WLM����ф4�n�_PU&�P.) �#��,�v�8���8���yek�k���x5Ԓd��-2c޺�����'^zC8V��i/ݻ�4|�z�|�&����vx[�M�ԫ1^���o΁��g��&&�Fh��>�� �i�#s���`����FA�Ž����T̀�}6�j��]j���/���6���Ҹݭ��]~���U6`83��ٞ��g�Z��mDE�k9�g�k��yR�bJ�.���󓌥{���"賿A2��QSC�;�U!�Cl���7zp�|����,���VӅ3F���*KKmX��U��&�R�!K��*�S뭍��s"nsC�^�I����F�Ԉ��+E��^�C�%��������N���̠�QMkEo �A�`�v���ԩ�}�ԝ�S��
����v��;�`�c]sz4�Ђ���lB�V�t -����܂�X�S�m�?�˂�qƜ�ٖrl#��ti���)������eH�ؖ�R�x[p��mhh��Rs��K6W���W��y�Ɯ�+|g���D���q�w�xnͤE�}mx�SC��V�O��inhcc�p2���D;��`ˊAq���%���f���cS ��F| ��� ͱ1�!�C�Ύ�1�/;��(����}u#dK�
��y�-1�[��\�+@���`�ľ�xt6`ǵ�$��ns�b��������5��y4��T��/>�4��傀�۲�'�]D���\�?B̻�/_��jm�1�>�}(���S�$�7x�g����]@�>}����^��hq�v��or%7�R�
!qYy����x �[����N~o�?�^����ٛ�Y-0e�POߞ�>�"�W{,�g��.�ug��ѢG���{��l:A	��7l!8�b��J�Y���{��D!rJs�q$��	) fpx��xy���D�q�nܖ�6:5yT��}Ei��RB����o�v�	�b���]8O%�.m[N�=ܠ���U4.Ma��g̰�̿�ݧ��F����g�4�ضm/���4�h���"O�_��D���u�HDM�ȭ�����]�J�TV��%b&|{9�K4o�(��`�� ��h��&#�~�ٴ]�;sqE�%L���:?�<�ҺU�.v�u�ǃ�#FjbJUp�\�K��U���ؓJ�h�
Ե���v��y���UY@�xVj2]��st��9��02���ϳ�4�D �cy$�
ECBn ��@�����������8̾���4�o�Ҹ���4[X�M�y��v�g з����}I�3��z���Q��/��9�'� �jɕ�[�ԛo��g��5�ǆ0��,��
��B��ÉQ������mPe�D/CصJ,�w�Λ\����o��bV��v`!�ora�U|�DV�����B�0�g5݀�)�`Y�$⥩F6��g�R�3ZvyO�@�Φ)��t�p�Nˬ�7��WS;�{�T��˰}�1�5Pk�b@����ݠ
��ì��|� م+��92*��b+O_VZx��]�153G�#8qv|�l�� �,�2aN����# �.�y��E�W�I��#�sx��D�5�vaݺ�H����Q��H,��>�O�ؚ���OX.���혾k�w�L�3@����0	��p||*�;��y$Y�E�!].�\���,fx�bKEK��"2?xn#(��-����ʍ�ã�3Rw�Й�#}��������iH���L�غ����W�ߚ�s�&��M��ֶQE���V���dA6��9���~�ʿ<e�EQZ�+ͭF�g�'���Q���u���k3P�Fŷ��xY���Z= �%7�G���˴W/x!�8��lu='�c�Z�h�m@w�����8ڝ����\g�����~-����}�ؼ���%ڕt`����'�~d���Q"� W���"R��vԠw����.��䈈i�u�`�%I��l��1�)�X�<U秅u�@�"�:�X��U&�fg0����VG;QGx��w�k4���3�9�!)�h�1�6��Y&4��?�ƍy�u�(�){?�wx=�����v?}�a��槈�}��㎜���-����r`����h������p�S�m��_L��1��&�D�:�R���{�]�D�����r;�E���'�HUԼU7�@���sh��X�8��\.���DN�Dt�P4�לA�&��L�'R��&_����%��<,,
Z\�b��\��._�[��j���B�\&e�=�L��&��)���E����QFh��X{׭��Pn���s��������Q�o��7N�%C�C�B�dy�<C/�=���s��[PE���[u��b^V���Q:�-��ok���ʹ<ю�zMȑw��[����"9������O���Q��V��9š��{91(w���1��>�����k��d)~w���D��0[���N�m����J�K/f�;�7�����H�rD�ɺQ�O�\��(��R}?�zb�*<OL�f�=�P����]�e�ڕ������Qv���0^��@y����f��5G�p<h�v�Y}�.�'��V����r���GAS��l�(�ODz����5��mSsq������w�֥nyC���Ns|a���K�?E�ϰѩ����-f�7!/�DH��9E&?�<v��l���0sB�x��~�6$�]�vs��f��esyXн�b���VbP���?ފ�����������?媢s�{&� �^z��V����裋i�%��a��*Y�E?�̖������+Ȍ��O���4fj����+F��^�Ts��X����C�T��C��aT`7��(��;��`.�S~�Z�poE���tݷunD��ӱ"w���ǂ�ȓ����Ei�bZ[���!�Z�/�цC�D�l�h��|�{��tS�IPH����?������ 	���8,2�#a��L������4ͭ)lX�t����R�|f��&A�W����k�����˃�1�[����"t����ߗ�����ޟ�W%d��YJ���ER��Ι9t�e3H����/r�eUjƁm1��$��N*�Y��p�.:�
c�7ťpLߧ��jQ���ZeV�,"t��ٮ��=e�/�-_)��n&_=��r ���TVJ��m�����*6�$p��5fw����] 5UT�ҙE4{1��w��F$����Ǘ�'_��:�
<VH���'k�eQp �qx!g����*�/ �!�6�6&H��_�3�[�P�3��K@Q����"Y�]p�L�e���u�\F��Q���-�[�e��{�cȔ���Y�|�E y�f��O3t!��A����ūB�u�C&�[���J+_*���H<\~~� ��@^d�ɿ5��G���xoL�TR	 s�=�LBf6�dq�$�9dE,)��n��N��r:�E��������٢�v�@x%��[�����~�����Q\���VE����ξG'Tl�+��4�|���9�(HpT������(���P~ M���-䜋��n��ݜ��SS�/���3�����ǠϨ����H����G��|p��¤/0�P$1I�=ɐ�:_���]�-;;�ܷ+i��%*��)�K�Gs��Ny7���=~��.īy�'�K�d3:�wr@��_��e]�g��Dm�mh�Ӕ��pK�����7��ׂA[�b������D���(?d�x��n$���H��$.��0��Z���2�Fh�߂'��Ʀ��U�r����qĞ_�'X�i�~e1>d����Ka���,;O[�>�e���?_�+i E��n�K�ZV˸�����=�����t���p�i��rRʹR?$*�%���@;�l� ��7��6��x��my�ul��G�=&�;]aSz�<^��d��	x�b"���obϐ���!<����Y���2}�����/�~�|����5/L7BHtD~X��h^}����/3Ib_�z���~���&�����Dw�:�Q;��9s"��xF�ӵn$���v�\l��zB�}%h�Ф����!�0eӔ�luMY�T�a�裉�\�p ���]S��h�.��K��"��ɖ�&��џ�*:!��n)s��?-�Ѿzb��E��4'姈�m�ϴw���u�[m�5�0��>I�^�=z�S'\ f��/�V�_��!qn�B�d̂�,G��>�U�ݳ��wWd�p�&cf�����݇ta�Ȋi|�����Zy�q~�t/�M��4֏��D�ܡlgP3#S�@Ƃ/����;�2� ���/=1u힅���Q�(��ά�:JV����G�
����KIc43��G�����,���6��Dpo!J��9����T[}h3K��-����j&a�T�";s���LS�7 6���ֵ��_x�o��~��P�d�R�׊�y�'9G�L�ᛟ�r��j�:�8�=�" ����fH��Q2V�@��������6`�/p�'�nQ�i�ʡǹ��n��M"x��{SXcܓ��3<�'؃ẗ5N�-AA��ujB�2���u�(��h�O?������D�"�F� S,��� Tkv�P���+�li�3�p��[�ǻ����!��31M}��[���pt�9Ϛ�j%o�t�o�{�p@#/&�ݝ�>¹=!V�b FL(ݜ���݅�ﾷzwgZ�9�kW ��A8ڤskbd��$���ɟ�A��Np����a��ψo���2���K��	�����L��� �d׋m����:����Q�Y����S	�3@�{E�$83s|��� T�>	��n���:I!׉��Y�5�#�j� �.Rv#dOq7~a{�v�Y�C<F@�;s#4>u	z�n�	����8�=�Ux�_%�237��wϿj_ؔ/���[�����P�i`�e�9KdObϼq�n�� ���S���6~n�`���W�T�N�˸7���s�?��0w��fO�7���Xֿ��v>Xq��
_>kZ��v�oأ��b���i�cTvVZ�͘m��_�KUߛc�=�N�$\Z4�<�����C�z��Ue�3Ce��S;x�fOZ������)�WU��޿9�<0�y4���hK��^&�O��8��`��2b3#�҉ƜG_o&���d�@�M(���*����)n������aJ�{j�_j(���i�H�LI��?R�k��S���u����U�~���y�Ŭw�ᖓ�b>X �'�V�1�I��{�������X�|#H{�5�ʧ�d��z���+�m���복ƦJI�����xmRJ� ��z�����/N�5�jf褷�r���� ��NvT��
p�O.��Vz	����#;z���H��;'��6��wg���Y��SlS��>Z��%7<��xJm�x,��@���ZD�Rbw�p�Ͱ�S�SR_=�ZH�s;x:HD���`Pϑkq�)lQ�W�"/-��dMJ|��eH��1��[sO�ӟ�(=zy�A����D�:=/�v�o�pP[,�Ք�9*ϭ���<��!��V2�[�����kH"��_�Yy��]�-��1�/����ϖi��f��/�M���4Z~Q^W��k�Tn�۞Oʥ���U׾�ش����Y�!��i�2W7�����̮j�5/=AwAL[�W��\y���y���J�MoKD}�9�+�����}�A����r>[	I���ln���ZYL�m9��ӐW�/}�0�w����Y���mt%�} 0!1��܍���u�x�$[�Rx-Cj�t�%a�zѹz�_�e@z 	�P���][��q�w���j�3���Xn[���t������+ tV�+�,{�bQ���Ǥ�����ζ3���³G�!�`�~z4+��}Qꮟ/N�Lq �eֆ'�!{~3�lO%��X�h����DP�����F���Mk���z��c*�Q��߉&�Ӛω�ǧ�4ɴ\8�`֙��cӐ�0�C��#	�n�|����7W6O��z�O���O}����j��Y���F�k��끏:O<:T�{��ػ����
��� �����owl��wl�/�Ծ��ߊ.�0��<Ϥ�{$X�*�2��+_M�bk���ύ
bIM�KP������Ϳ��,q=��>�e�!6��7[�c`�8���f)
u��f��Np��M1e�9t�8�L�}(��]�T�$F+#o� h%��Ȑ�yI>nF*L�^ͤ�[?�7G��N�.>�d_�<D�`s��R	q1��vm�(1&}r�実��~%RkK(�	�b���j�2ѭ�
�H��)�FQ�>ZA�,C4#Qb�No�nU��p1�ҿ��̮���7��&�G<=��5�[V����[8�����:���Z���t��!��Kd�s��j_�V|Ʊ7�J�[س��`��Q�쀠�<0�Y�i��-�/mʹ���5�����^��0dǝX�����	�7v���*���ob,D_����/E�u���z/!)�ܑ��Pi��p]'���⏂$�t��v�b�5/��z7b�Snfoh�uO�s^��)��;�ؔ��o����C��S}%���O��J�iW���p+��̳��	�佚v"+�W!�$[���e]kF��z�[���~�f!��.ň��~��Gި���A���6�b������+�X^������B�;���M|L���8r������8 *�o�3�q����^�'�2�W�B׺��"y[�aZ��D����s�D�� �Tu4����L:sP���!���^%a��x��b��ǆ7t���'�IV��.4����P��'\^��Un�����10º}��N7�9=�5�:q.��8���.�j���W-ca�R��;+ɢ����.;LR�`�z;/3B���";����!�l�et��g�Q���cp�r�2��F_E��Ww�A�Y�_\�lG~h�����#8(L
���|�NBB�㻗E��zۛ�6/��~��pW�Wm�2"��Y��).#�z�?�8ToMn���'���I�  ^��ƆG�c����b�o��e{�����x6�N���k��R��u��
����CޫM��2$�t����d�ݹC�l5����rR�es�eL8�;���j���Zr9
ڭ@������Ǉ�:���wӎ���1�e��I��#������.ǽ�7�
,}7�P4z���l=��܎%�-'�i�^<�
K ~>=0�� +�J��Fq�b�It���|�0�V^:�2���1�/���6��j �z��ή�a\�2Q���~e#oXs*&�4�S{��4���CG.e�H��?���ߚ��	)�K'|��3�쿼���)�������g�[EUCe�����4'��?ǲ�w�z��:�H�G��c��E����`t�go�yD�1E���jJ��m�$��'�>{m�(D��bY�%�bT�c�
3�81�/XT��F�j�oL}UT�&�I�$��Iڹ �C^s%_�Tj�mp�8���'Z�4q9�"nj�.��G����b�Q"�s �v��1�-��������|kB�|q�	m\�\D�#���
Q���T���N��ax��T�����*bo䋇��z��3�	������`t�ɲnh�o�ʡ6�ۊVЀ�[!~c�d#�� ��f<a޺���|Tj���n�������}l?��E�������h؏�fJ	Z`���]�l�m��m���ͣ]�5<5R`<IWW�*D��0(3��; ��uv�\�ohb�0��L����3
����]/	;��߭X���h�n϶j�H6y???������n�O� � o9J�?�c��i�M,�����r���Q�N���������.>�
��#�|*�P.=?�)���[e���Y�o�?�}E�#��?�_�}��"��"��!g�c��|��,^��&���r��w�g�"�����G�b�A&G���w}
�G*d6����h� \g!q棽���H 9���J��v� \1�����<k�nC�>��K<���t����u�x�@1Jr���Ƿ���gN'��W��J�},F�y=�Q��v�;22�HX�S�����=Jj��%#������G���P?�ɂ �3����.V9�����T���uE���F�/���sα��T�*L��#���z������/�U� ��B���m=r�0Uڋ��_�O���ى<��PQV����ڪY��Q�T���/��e�~��]kQ�_�B�D2�\�B<5�oiW �-UKW��-�~��=XX� ��T>.�bQ�����r�+��]Ȭ���-���_�� .��5Pr=����$���-�V�A�o)EڌQ	Ĭ1kdR����~�&�q5ҏ���Z]]FɌV�oE��7/�_�"�O�<6]T����
؉o��g ؖ��3<R?�Wd�p�mI�ߝ~��]����\��=6DZ��鈾���%Xo#��)���J��l�2n�̗ܵ���u)�c�SVE˶=�����ہu:z��f�.b�����-Ў��?����΁�ힷxU����)6�&�)qm�s�͝�h�di'�7(�y�݈�;��N�N,�(mp�È�]�j��)OGgt ����=6(-� �����*o���S~jIi���'�w�<�m�i2pj��s�P2+ИVu�uh����>Aڦ�y8o�� �� L�qw�޺�_ ���`�r#����NT�.���Yu����������!.z6'a��K���O%5Q�%a���Tr� .���QrRM�P³��Q��ցg>�ʾ�b�"�D��X�%�d.�l�RO!��۞ir�W8���=V�/��(7��i���6x1P�Ѣ>d͟�]$���v$�Y�fy;C��@�ٳ���Ka�>}?������
'�hS��D#�wn�'�~$U�����e-��w���m|��ev�`���@ڷ�ͪgH-bH-��+�a��bg�q]�����ى}$RtQ�}��C�T�=����J����h��z63��'���s�¢R��J���)�$}i�,��;|��Y8���22V-�^5։��mAds�=�/uG'�*�)%���4�]b��& ��E�<�}*T#�LaaTN��_t��k�ݰ�/��u5�(�������N����,��0%�P�ښ�$rLt�af�R)~��r�{E�y��]�����(ѧ'kҶ�":���a���sy�F�OwG�w|�)�@�T��Oho�x����Fݢ�-����5��y�<�>|ͯR�}����*�L��l��`~����v�b4��p��&���1斃j�2x���c�R\^�J�-�T$'���f�b��w?�/��Y���p�Y�2n]2yދ�֮��'Ym����ӫX�&8ŵn��A�������:G�ز�j����$�B�m�ˎ����+벢t~>�XP�<�� McM�'�F�ʽ0�hQ�uci"1N���qrZ�'N�z'�$��=nI�f*���8���	�!!`NE�*G�/���͕��f����0׵̛/�!��L�qN����#�,Y�/C>|*5P��-(�X2�r,���%��lՑC���ٿ1mr 
Vj��ӧ�H_�fmF#�P�k\�u!��|5K;-��ܼQ7j/��4a+x��t��X~��3kI�TӳT2��Q9(-����t�Ls���1CbEX;e��Г1ҧ�<�e���K�����P[��\���b��Fk�e Eol\��XXY�2By��$K��,sʶS�Ĥ\��ݱ���Y��Y�������bA��?��:��$��a�ּ�!�DbcV���~����Zf�\_�TW�\����S�W�na�]ʓ�b��-�D~6[��9�.�����n~�@��G>!-q�����V�|oW;���	��a_P��bc�Y�d[F��У�b�8�� F�՜�q>���9N=�ke�}ĸj}�P��g]�l�ݼ956�A6������V�tUN��&��|�$9`�(�;��V��PY݇Y��� 5�w�}s�RQ���	f/ ��1f-7y.���V~ʾʟ�\�n�{�u�U:��lD� 1ޓ�� �l	���[��38E]�O089�jԵ^��]��oIsx@��w�}����X��ŷɂ�Q����,uN"��/��鹟�ۈ��# �mF�.to�T��|�zo�G�%B㳜F�~�s}F�8(P�����p-�����&����n�[�к�[�B�8T�_�z�>��;��ƿ~��Uu�W�(��PAx�L,�����z�C���q��:L�E��9>J�n}���$.������ej����՗��po6a_¿k���kj�/�WPGr�S��:5;���������f�%�#�E&g(h��}-8[��Ă{e����kb��C���ݝ�rmd?�I�	�B��p��zf>C��5Ie��*�V0=��p������t���
W;?��D-��2'/�)�Ȧ����L���Q�1�&-⾜�ԇ��q�(B����1s��+�j��i�Z���y;S��m���
o�N��A�S8��_�WcI6�B�zj~������f�ɮ/�ZzLɩ�LQ�(��l�R\���|j�,��;իK�
��@K��:(7�Z*��C:8��4�̣tY�]���uFN�p0�d]J��#?_*W�;�f���m�nRkx߬��x�Q�d���@����ɤ�7I��ݑq��};F.�
���[&l�閧����>#�`�n�#5�$���K|""4÷�wx&888�777���-����
����>����ă��'���k����Z����9Wk ��-i��6��c��K4���ܖ�K���d��Xb7|����l=Lqf*l�s�
ط�ܼ�NweY�/#�c���^�wv�:����HrhJ��Y���(���~�s�-�(Ҡg��x�.�HO�5?SlJG�@Ŷ���,K��S�~B~�e�`ϵ�oG��L�H9	>^��o'e��B7e|hz��o��(��b��N���D�@��v=)N�;n�lծ�L���81J���O�hb-)GuD~��nO�����V��o'b���E��3�V��)n��KKw�O�{��i���\��(����ULp t����<�J_�,z���~�5���yOZ�OG��ѯ�
\E���Uht��V����
摃�]�ł�W�ԫ�I�)'��C�mx��p{������y�[�*w1�Q�dQL�4�i9�+e]5·�Sz	�"2�,��/x�8�Ŝ��$nT��
�A;]n�H^��ЭQq�`�	������f��-#ae�T�d�32*�f?��>-�C��x�����dR+�����e�t��)�;'�2��NuY���;a襚���#���a�9��'̛m}:�X�Uy�y�W{�Z�ŧ��
^C�I�e�2�:�� �=�K%,���5E��H�K��3H0�'-�+��!XY�iV��?�u*b]��p1M���(�S���1����s�79͉`��/1��%J�r�Sh��kGJ��<1��hcG[]���k2�+��0������ʇ���˺O8���'}	U)>�l79H���xU���+XG`=1��ל?��w���u!���G�Y��c�./o�(�;j��{E|[7��+$6�a�� ��eK׺�"��M�"��EeFb��*�'mL*l��/�K��C�[7�;A*7�cTD���� EE�3��O�?��=|�o��-���q�Qt|��j��-d�%'�1�"�5�4��gJ_����O�p�y�<L����z1ܦs1�����f�^�σ�)��+,T�:j�*jq���҃IwK�ɭ5�@G�v�4.�H5��O:G��T&���g>Qg���Z�\'b:����@@��fD��6&��zk���bY�O�	�	����A0U��K�YL�}n���\=-�����%�w0�bG��&?)������j�U=UT2�lS$�Z"�(� �xR�.O��R|��60K>�⦰�+2����~e.!�qpG��.�S]H>k�i#��䞽��fx\�zn���X�a)>l
_�P}Z�W�Rǃ9�W���RRߍ��'y�GiV��ʚ/����3#��}	�n��7c�ZY����u#�S��?�{u���v���ח_��6ے���Df}��-�F�J������[��%�#B�GDNl��
�uYfMe*���Z�U���L�p~Km- ��٥�"r�</��b�tgQ)>fL��mE��@���Du��u��5\U�u��y;b�oCc�F_����{��m���K��7�Q/ �'`��t�W�����:X>�-���_�V�f�������O�RN��"�5�"�����˒�ڧ߳�e��K���~�l5�z!X�Ć��ВRBl@�Y��M���תP|O���������Yօ�����Cpw��Y�!www'	����m}��o߳�s2������Y]�T�SsVw�j4�{��LJ�0�G[
�)�Zi��g1�N�i�#���:�x����!����W�a씬���z�y�]Jc�]!���~�$�3��/d��z?h~����q��?�L4���^�c�<�c�Vt�X�д�7�w至�S
׳��O�Y;ԩZr��sv׹9�h�kN��h�"=�z3f�vܠ�7�V��L�{R1���3�T�t�f�8��â��|�~��%�1��fg\���c�l��6����<9,�,�oG�&�l�u��ڷU����������ƽlB��݉��_{���K�Cm��$cj��M�0�qwF����oL4�"��;]�����%'����>��`�6��	VNb���Ā���MpK�Q���4^l1��V$DW$$�����'�"$J��_��Y��]�[��|M'Im���1�<�.?�D�/��HvZ"<g�� :�fE����-r�:��ϲe2%ȏ��m��t��q4�>��w���,�mL`��P�����5T���$��|��zb����!�6�e"��~�JU�р����i:uD��^��C|���xX�^M鬇��t�|{�4�)z�^����ZX�s@����>pt5���%J���SLh����7����܈�K��2�}{�^;��F���V)w����¥y�T����t���)su�	�D����B�V�P|���v��'��x�p �B[�V��}�RN(y+n�'�;U�g� �F��J"$K��ܰ��$�C�sJH�e����%���T}٠���I�3�o�h�����/�~��P�H������A5XY��tOƇݍ�a%���@��q���qN���Wi4��2����:QW�0
�c�u2��s��z~����B|�@�K����C�2[� ����خ�� ����s�%���P$h/�ޤ<.}S�|[ �^����/Q��N.� ��ړ�	|L{R#��S��݃�Z�I3��]�t&[ڜ�[���:��h딀0�}����l�}T�a%��R��JD�M��c�i!T���1�|�Ce��M���:�p��� I��{Eİ<��$�؅�$���A���(�P6�duR��?P8H{p�zb6e���vF�V��������/���^L|Py+�)����>	B��͈U< � ����9~�A�������G�>�;Iߵa_��.5"H�=BI.���Qb��EOD�N 0�#M���K�U��"D�O}�&1���\��a��k���$9ˬ-��<AHʤ/��
C�nH���5+���������!����5��^���mW]і��t�z�m%$�Uނuٲ�����":xŹy�33 ��/�5.]�:\�v�,ȳ`��z���a�ZNH�씒Z*�n|�n��:��,R�<G�?Kc=���L��w@ƪ�^ؐf�:��b���{���*v�$�>��	����+t��om�m]�KpLZ��n����t��<�Ä�ӣ��$j�s���'~[ˇnc� ��B�{^�.�u	��뜮n^y#��͝|��f����_@�v�s����4z���� ���<&wu�^���H��a ��ި��E��`sKa��}���G��~�.&rz�l!m/�#���6������ I��.�<=8x����/��)����Rպ�+�v�k�:��ġ�x��[��]�o_V���ؾB��C+NHD�w�%Y�С�)�ن���O!�ߵh7�i��Qx�x�׎��;�T\���A�"Zb����*=HX<��gB�0@c���5��,C]�����E��kD��1Z^�d-�_�,�G�ѝg��1ڱ�X{��+]�j�P�e-yZ���[je�HB'��i���ᤐL��xИ�zv!�}��e��H�ǟ��|]n�G�=�^��&��*�,@h~Lso�<��.,1�=)*�v�� *�1-4wL�[�;�t�I�������� ��;l���%Y.
-l?��C�6�܃�vC��KH�C�^��8巰}���.���ӫ]�K9�q6R�D����%]g����6O{��_��,b~9���N�����C>�?\��>������-��%%>.q�����q$�e��]�����U|&&L��$�}����"��u���v��b�R���%U�����.��+)��2AE�j>���u�4�-o�|�_rr7?f�M���$���0u3�����p��]�4�=A��'�V��_V�K�J)��\���������d�ja,b<�P��FMɻ��`MS��n��=���N� m��k��pD���K����"���P��t��5V���n�(f·��<nit�<�~�b��ӯ6��mt;  �]�V!݌ۛ�f���N�[k�( "yo��_�;=UQR�9ل�3��z���{}�Q�l~Y[ԥ�C31���|�`�\;JG���"K�{ψ�C������9������3��O%���t�)Vi3�#@|��R(Wk��vJҎC�J�v�E��F��'�����iX������a�ij��Nl�-�k��N�� E{<��O����/\ļ3��T�˖lHқ�+�i2��!	�7���4�׍���"̡"�5ж�0�?1��Tf�ģ���Y���4�5S�H�,�Ξ/���hS�ab�E���	�J5F��Ag���w>Hu�
�?�-�ߘ�=�
ӱ���z��Q�e�%K���F�9��y{�@D�����md<Dy�g��l��ba��#���[�V���(�7Y�A�����k�S��Ľ�)�Б�k�S�ZƧ0/��θ�N#�Q����f�/�?L6D^.?���@�'���Z��a���N4����(݇����_�fu�:6/�Gim�<��(����J^����|����^�B\�����/rdj��/�:L3ܹz����?���U�t��GYyg����i���J��ٲm�����������!�E����M�Slғ7d������*�7G��a�t��{#���Z7�,��w��Zj�t�d��#�:(�ZV���i4!�JVܷ�y�W-(���f�+w�.�g�#R�As�9����뵐����<�?fi��hi�jtӬ�}�XX�|���������'iX�}�I�	�lX�+��;�Q�U5�A;����xC]�r���&\ޫ��Ö�ˆ���'Y�k�ۀ��d��!w�����H��u*c�����O��S�0��v�t�]��n���ZӲ�AT��X�]��,|��LT�b���눃���|�{Vy���5[�������!����+�kM!x�#ٕ�L�{/G���O�h4�0ݪr������j�<��]
�o����R8�n����tX�a���J&wi���f>����r\�S�Uo�l��R.�,�}�w�i|i��1�V3�x[�/ͯ�L{	�K�fR�y��1h�"&�Rb�oH�$�>�&o����� ��zf��'!]v�S#��)�A���3:�_����j���
�0�����\"�h3K���_:Rݭ������?����:��ٕ�5'�ҧ��}�:P<;ލB���b!�->�p�U�+�-!��c�.T���dS���|2�z��k�O�Du��!�!�rK��Ԡ�WM� *I^��Z�����S����9�-,I��<�e?i�$�Ϊ,+)��Ǐ�kӷGנ�-N�W� ��ܴ�{0j�z�Vn^�W���j(}V_�o���ʊPTꤽ=-���al@氯7�;�!������N����z������FP{�Ѿ]]+�wZH��D��,��_�i���b�!�e#p��}���q���X�ƨ��ud롢u�������QZ(,͹���O��F��4#��A2�f��������<����yvt����y	��u��$�s����es�'Ǜo�[U3m���V�/^��^t�
���!�$���l���P����5X/�jl��mm����y���r�0�{>б'`���O�R���:p���������M�w,KJ�~z��mۭЌ�u��ظ=��N���} �B��y��RU�uS����ڝ\v79@?ܓ�n��Z���f��o���h��O�A�g����W��֭FmF�������El)�3�yT�- �n(��#��Xr.-x�R��Z��4��>��<�CU��5���SY����y��8�"��L��"�o10�v��<������� n�Y>�L��sI��6��4�mCA7P���ZU8�،�Ȕ7�M��<3|8�h-��i������N��W��8yݯ�]�P�L��bPچ����~͟a���F���Q����@��D5�����uT�{�abXS-�'Ŏ-[6�ހ`�q�pR��޴V�����#�m@EgJ�M���"����.X��,~��2Z�2��"*tv�����Ǚm���c��O,C|o9s�C��S�F��G.*��9<L8���:<��k�ֈϵ�.рP�^�f�$��l�	o�	����bT�C�T�`�
����#�n�EB�Oll�{���xdێ	y��1?�R��7��uuǰ)[/�_�x�	}b砐�uJK����Feb2]pǦ��<~�O!W�Ϙ��XӺ �J�7r��h�b�O�,��B\j�"���M�K�p�B�+��ϢA)��TɊ8I{lv��� $��*�dȸ����ō��ߨ��<�ر��Y6h�&���-��\�*�
��UV��u���L�sH��Nq4>��A}=��4����<pupA���	�4�;z��ڈq���Q^�]��,�N@I\��g��0⺫p�H�ڟ5��<`("�f]qØ1,1��e���,��1z�H��'�t݌%Q�ԈI������S��e[Zȣ�|9�,��H�-�����7[�QT��j�P0��,ZZ�2"�q�����#�^�G�u�%5��3y�f�i
����i�t�߸lތ/��4��f�%DJE��hJ^wy]���Ѳ��#	fn�Z���$��Um�Ł{'�ج��׹���2��#��9Xk���V���p8ȿ�AV�Ծ�a�	�#�h(ߝ^����K��y�9�$����Q�X^�pV�ٟL�he4�v(&D7� �(����+,�e�a Å#ƮB�c�N�A��ɯN��T��Mv��RP�.�9��v~�sJE�����+mB�
���3x�G��Ӑ�M��ՍB��I9�)�f/X臬�jU̞�f)Ǹ	>z��/
�E�,�k����ѤԢ����uM�g��:�4J��O�&��m>�s���m�ҿB>�'�ja~WDy��WP��%�|;��5֔���R);�[k��>F &ƣ'@����?���DRg_�i~b��a�u�fl�8��kp'�c���6�{���HF��^u����C>�	���1h8�9�|�����q>��yvS����i ����l�>���[�$�
��rll�G��
95��MTDb�����XYQ�R&e�2��bL���F9T�+�r���'{�=�FI/fF}�b
��I߬:FRe���T����\�rD/~������^��#@�'�.C_�LAh�B!�c�حk��g��[/J�}���B��*�7��jRmz���.����f&"�46�7
����EE��Cm��*�U�X����<�Σ�8u��1��Jgw��7�'㷁��;ӿ�_Q�W	:��f�2g�.J�\�����׎�:o�#�/Ԟ���.So�0����C�}fj*x~~����޴0�wy"��wt�m�G��Bd����T���7Gji}�W>��q�y�:�4ݢ� ײ�w�|�������0^&�	ʅ��>�ʥ�U�B�#b����@L��U��C0�h,��Ư���/E[¿S)nw�fz�[��[�v�g<H�s���bi�΋�Ƞ���3��q�F��v�֖�"M��	I�Ю���bݞd
xK�����+��E]v/��v`_I��H}�z�f��>@��6m�����#ڰ����*fJ�4�	�DB@�4���T&b�p%�~�����%VDp��'���ɯ�d��V�Γ`yAue�������-�3#��F�	7�p�����D�y��WG��ja��|�Ҕ�y�����w9��Ӯ5����r�t���b�*�X�L]j$#3XQ�bU�o���xC1fO��?NР��@��v>4;kR��\�ˮIw�4��f��l�����ǀHÆȈ����k��y���
��u����Uw���X�<[��;"��}Q�bO�p�PW�'��m����^76�3tpB
��o�n;ÔZ#v�#Mn���
����>sD��HqT��G��m������eD��Y�Oo*�͊/R�uW�h<����t�/�������l�!Қ�ua|�i'�ɑ��q�)l��Rk�����=ٍ�4�8:B���9BU��g/Q�(.�|x\�b�}�Q&NJl�S����g��&������XC���8;����s�.��}�"H�sJ|�s�g9.����A�%+��I�Ŏ<X�|@���'b;���������/�ykAE�*�&!}jf*��l��
#&�����S�7d����"��:�K��?�5�2ѐv�� ��޿�s��(
�x��Z����p'��n�"v)��)	9t�9��W�hD*��%�X�w���YB� S݄�K��N8�&�,���T��?��ߙµB��i|�=-z��G�ST-�P�b��K^��.~��.t����ݽR�����Q��Y<lʠ]7 ��4����(�{��淐�����`-l4��=�*1]0|SNIm�ޔx��Z�%��Ig�_9���|�(�N���a�|	g"�lF�󁝸��u�mEBk��6 �86�a�Ca��ɩ�3[�BEaB+���� M��п�H���a��H>ЕS�;��jp���?+�֥w��,�-f�b@W��!�:��� ��%@s��	X�?i���5�E�Sa�+9��-�S���-ҟ>���X�뽁݁�lQ[�bɭ�!��罛�o�������д��	�>>�Sf~҄D���ⴓCc(�n2����kT���_�("zֳ�����V4/o���yٻ�������7=��	���Ss���i��E�X��#��i,�!bt�(����SZ9�m~c����'�Y���q�j�QZ�H���q�sC��М�4ϑ�ww)�����2��ڠk:v*�sM�������p#B��Jl��L�����mZTL{��(B�`ۭ�" [��L<h,�>Fj�1��xw\�{V߰���o��G�B
���w�-y�Q�I��2��*��LA ��쨨�$�C���}�m��zX�|p<��v��A�zh�E?�������ݳ�I~���p�iM⨨�fGA5p̭kR:X�Q���,p7r[��#�Q-�L�bc`�Qj0�<�h;�G<�T���(���aa2���)�
z{}�ti{�t��x�h�������5m��z2�t��1R�"r� ���I?\�я�s�P�� ^��.u8��x�u�l�
���t�:���7��%iwQ�B@�bC(�:?s
�� #L��  �&��T"�k��Y"�D�vzs��&q�M.�=��b<f�����P$\�����>0[sZ�fȬĆ��_�kG�ɇ�_�a���'�<�O{�m����7����E��G���=�̰,�@߲d�T�p�fg����s�<c��M�l]��L<:�}k\���������֏���~�'	sz�{�K���҃�W���v$b��7��߁h	�<�!$�H}*�H���,�%{�<c��tO[�t	���5�����Ǚ��_�I�~	��ތ.F�Ӄ����$ٜN��@pM}���	���c���ݟ�޾V']U���JٯKOT����0��!&S@�MIM�iwظI��?f%�F��l��!�s�l�.oϣ�㿴�3}c��()��VռMB-I���s��<,�}���Z�H<ϣ�4u-<;>�@U�����u�^�yą&Ox��븞����z	u����C�1D���$N Ø+����n^�RLbշ,b�p���z+ ��̡>a�f\��s��yF�����?�?�-dI.��	�T�F�VV=��q��"�Y�R�v�m�R�RͿ����3���P�N@����u&��t���X���~y�[c��Q�cp!c t�4z��Q=���-��2��5vsJ��	s}��N뺰�5�hq�J�|�1�"�a6�8l���_��������ι�j�P[��x��g.hl�"6�������c��O�@�KVx1s������;�z�@�1��@��W�	�܏�#6���ZRkf+칸
�r=����2��\}~��L׷��&��(V�I�Z[[g&��������1PJu'a��P�0��k��y�p��L|���	\���!/����(����������O�Πu���,ϙ|d�9��RM�c����ȁ2!j݉ȇ�_յ͕��B_e������]��ҥ�K��kl`e���G3�E�B�"J�<e^O�(e�0�| ���1�N�[mqU�@�`$6p8R`�����6��M���b˳¬��/�{C����J�w~�k�g"q<e��I���F���9�.&� K�w��M�1b`�Xo�Pw�J�~lUԧLE�|�ap��S�H��IC�d>�Xw�����H��E�@�����<%c;o���(����3+k0�^�2좻�f�s��?�.�KS��&�W�o���W&�$\|�GbjQh����ԀY��d��+TDkmQ��q�^�\��G�U�3��D��_@d�n��e���������X3&��Q��D��x��[��f��� �Q� ��Z�� d��C�i[���������QN��l�����7t�	m4�Ӻ3��Y�gg�ry�J�!�S8l]2�+�0�p �L�z�����I�Js7�"I��]yg�NIP�;$L�M�VX�����]�n�^�ueJ҃v����zg�K��{���SɘcE�`��vw�8�o���<R�=1�^���f�=}�m.77W�GlffvF�h>]�&66������"a��[Ss�xq��,��ϐ|fV���Z��Z����|~�.#��z>�v�O����c,[�1&���Uo�D�;��Nr��vV�3���.��W,{.�n��&S��2��3��$��:��6z�c����jE�#c���@��~����L ~�!810r ��3�]XT�DV��v76*!��W#�VPW�s�z1���|��Z9����d�$w{`4�e��_c�p�]�m�Q��fu"燨�����Y�@ +�H�a�8�O��!���!*�ӳ�G�	�k�P�\asm���.ؖ�or����8��1`IN��7�8�r�T7��з�3j�� ����"�	�����u4���f#����bs�����y�u Ona)C�ϔX���F�0箹B�g
�li>��& ��f�us�t����/}*X0[�"@NI#d*�?�n�1����k�o��Å�nN��(@	�����w" 4`��x�i{��݂�.f� �7��n���D!���_2�̔n�)'��v�/ՄZ"�<��z{����˩�8�i9�L��A*��?湊C^Ԩ�\ߗ�_j�6����j_�D�vu����C�ˤ���Q��l_^^6_4
읜�҆���d��:�>���5��p�dtjmK`n�n+�P6٩n.�hbW�,����O���ƵS�d�tl��ܪ�Z.��SR�b�WIw|�,�b	�K�������;�0]��O���]���5��<�I敨���H�ϐ 7&R�-P�Ҏ��?󯔤4�)23��9w'] �7uVi��uu�U^�- PNM��2�7�Z1�j�ڭ�Q�w��Fx�#(Ä �� �[�>���|3f`{J)�@_���\�Va�t}���J�RQ���*�!K�s�x��e����x�� JO�}KIEB��s��ü�{e�3"��#��H�m���ۉ�H���~r0�- �g,Ӎ𴒦?���/���G�?�Q��*�ww���ca�@,��6i��yh�Tnߐ	
�S_CJ�=3uw�|S
��zm�#� ���SVd4L�hvV ��Z�ʪ�vo��CmP��}c���Î����y̧Nse�� �&��� �߳��^��_;�9�O�q���z���d�S{��Tֹ��WCעi�C+F�$�x�w=&�Iɬ5�O��j��Sq�]�ӽN���0��oF���-~�.)�R�=%rɄ�R�#������3�$���y����P�^H����ʱȑ�D�,,,�_>�}�V��b�E}�H���z����t��n�Y�5�x8U�_ƶ<�#��.��
X�-%'�>8���p�M�X/˷����r��mH��B��]���3������B�P����z��{��,��*�|��w:���Y��2��S)F������jR�	��f�]5Q���@ ��������'M=�6/; TO}��&��\oY�v�)����g�H>z(ǯ�d.GU�U࡛�f+Q̅�P��(�&���S:F��vMڦ�m:� �ٔ�jޱ�P��*�lK��z�f�n����_�㨨0b� �>�����-���5�v��;iI���lxp�4Y�<}��Ns7�����u���N-�4�'knĬl�t��	g4;k��ٺz�����qPŰ��	�	FM*,�Tk�nY�F��a����>�o�p�F������,�F*ja-�ICJ�TDF�)ȡ�3�)�fX;����(�=�!�ܢ �M+�at�U5ڒ"��j-��� ��>�2��V�����S�v�6��c?�QW�Ęe'{ә:�؈`B�4tg�e��o�������OZ?A5]�W.s�A�-?�鋚^���oo���6���X)ٿ�r�o��~Q� ~Z��JH�:���>}������1�11w lni�z'}�)"���`��K��_��(�'a9)^�Sk7�r���#O�%K�X����k�[O�zt��xd뵹,��R���E_��ʲ�V^����`���B�����[�͉w.s$Qq�n|�Mb����0�ip�MHP`s<�
��n������ވ��n#>+L�;T�k5;��]��Q�,����5�+KH0������X<hm�J�,��j�NN[�r��N���Xd���-λ�>ZżWĉ��Yץ�ɝ�pL���GvE)z�G�H�:FGm����	!�E��LV���D:��Pf.�v@�|R�d�^�8
'�u9���Fĝ��?۔N�	)��L0�%֙t�-�`�uםc�ٱpdN��և�3��0vP��0�u��G!/�0����턝fA!%��M���/�7��
��&	)10���U[�E����ȗW2s8ɢ�r�����e8�%�b�cb���/�j��S�f)�����ȝ�X#�;9�g"bfe��T��$�2�CZ�I�Q6�����!U^�&~����|�2�����=�pu9�����^o�L'}R��8�u�bN�q��)Ǿ=Т����'6^�z�MQrBJ�M����G�2&���\��h�������nrT�F����x�RGF��L�H���{��E9Z�t��W/�,̣_�L�ݺG�|���z���}E2p9K��x�D�/0WY�0֖f_�ݼ����4�&,6����VWw��o����y�>��:�{��foOY`�?�GƝi )�3��j�k��bEљ�p^��צ��on}�ǎ=FF�ƃ���6�@�TW��^��M�t���)�k�܁$�i{�̄m�ƒ�����o���3�%�}}xx���`�����/2qe�);)K�RW�W�Ia�5�����ja4��;�dg�g�ݒ|-���Gʆ�ė�Oߔ����>Rt(Yк�nM�Fx�ϴK�}�<6�����3������2���T�ښ�Q[9]oo�jMk�|�h}�H�V,�8���;4 `��x3_�h�#�v�~	�C<��+�x�/�`�HT�
�I�}�)!<ĩ7 �퇯�0����<!�T�L�L���r��>���wa����T�!�^��Rg8Uj� �v�v),�eK^!��J�c>�q���v]��S�9�a:U3��H�[w�c�h5S)^��yD�M��L�iRO]d���'�71L�n�bb^g�|g#�+��K�Ƿ��nM�-���S��U��k�:��mʚ�^g�#��w���f��Pu��}\���\�(6�����m��HV���y-@n b|K`���*�U�ſ������뛕ٜ��XUTP�{U[V.w��5�ijޣUY���5���j�m'g,�n��Cw��&���k�x~��X�@�DBr
��82\yh./�.�i5�,���:i�2�S�`X7�CJ�+B�	��F�w�V>�+`<�#^?�Z�����G��kϒ�%K�zc��1&��8��_i	�O��.�͍k����-Wr�ì�<wN��׏�����:������=DEEŭ��R��I4��x_f~Q!<f��r&�߂��HɅ�n��R��@���xS��T�p~�d���x��ym��AN<�c������Y����[�/Ķ���m�4J��@3''ը�{��� |/��������o��`�פ{�Mл��.⽥r��Z	Ks=n����↪Ι�P:n�t��@f���t�tJ՞ǢvoX�̽�Rb�/J�,J����F="�2h����v0�EQ�����ɖ[X]]%�}�*,+c2`��h�:<<����Y8:x�=������,�}[�d,��X6U�zk���+g7��R���lI	���-Wh۩p�ڠ�3�9���8e��S�\O:靈������ׯ��_k�p�?��&Y�T���T[�]�c��ӗ�r�Q�8��_�a�<瓯�D�x�ژ��ۮ������N^/?�<���!�.^U����I�d��p9���Q�G�%=dz���4)*#�����=��8;�R��	6��1~�}ޞ�7�N��@�a�g�ݑ�Qi��x�6=��ʜ��<�+k�ںמN��<��;c���t�r�k�]�>��COS�#�V�A�3*��^��GTW�5uʓ�4���>���y��q��a�uc����*����U{?��5,�f� ˰��Y)��y]�mͭ6�L,�֫o��f���Po�ff{����+<%�}:�9(4Y^ 1� �����NrW���%�}L�)�p��<6��{���ld�cݻS�ب~a�	���"����K��}�\Wee�Ur>ٟ��ՠ������G��;���k����\q�S�S����1�徬�0:�[\����*8�Il��I_�x��@rr�ǟmat���a<lV�D�d9��:ZU��s�F!�e=u������2A���_t���tM��B�K��dmfZf�J𸸸�ֳ�z���p�i^�����rW~w�u����f����z�z7h#��[�:?zw���j�s�61%�����1����u3K�2�����`�(Ɉ��>���/ż�o��ҿ��!2��)�-xd5AH���ʲ�0��Η<&��A���+�&o�'�zz$2�ǯ�}�v�q
�o�o��t֨No= 
��)�fШ)̣��X�j���
��W�1F����Bag���
E@�0�㢔��ѭ��15��̽��8e^x>�������킥Rv}9�����J�Tx����}��������	��-��ۙ�>�uW�k���n�c222ǦC�$
]��򚩆�V��%�z��̰|S��| �V��JAO�/����v�|Q�-��mx�2��ׄ �  ����I/�=��"�*_���@��,(
^|u{0��nP/�����v�x�2W�2���N(�4�R��[��p�┉�v��_�D9���I���{&!����<�K�'��`q0g�H���P{Z-��������`�(J@Df�T���ג���&&R���8��חӳ���@�Γ�D���R��������&S҃����(�hN������|�z���|v��k&mI'W�JS,p�P�Љ��_�:o=�ٵ�E%N���n�����o<ކ�"�[�Cmm�QF�վ�@" ������g��Tg�blc�i�gWZH����w�efN������/ Ұ��QϾ�����O/ӎ��l�p�_OT}��f��ogI|�	1f�t���~�k�㭤��(�xyyid��abq����9��yg�>��o&v�\�;-�zM��Ʊ
�&��`7�=ʑ�k"�>��#��emJ���r��y޸ ������x��d^��.���ԠCC��D��[�Jy#�1{{fc/pZ�_2�dH}@w۹� `d�������l�Qx�Gr�3j�R!�.�c��k^CIm���T�ݪ��%!�M���x�55c��e��:h��-�L��Vq0�kj6 ��d�Hc$���w��ٰ��d1�atk��錡u�{	I�i� ��Gg>�rNbB
sdB�:�w�IU^�^̪]��������;��r#�c�*��(��k�7?��Hd/�F��?�dQQ�g}}�$��'1�"2��$�����mZz� )��h�4�����1ǳ�v�A�@����\����:�-���.�)�g��ƷNh��u樏�Axv��G�x���d��
��/�)��&Cp>.ܴ���[�]G�Ϳl\8�E~637��:v�܁�M@������}FzU��h�Y��s�r� #<4Ku���!�}[�����ǳ�dx��o�B��M�˷L��o�Re��m���󵒴:-;WV�O�A��Y�߿���=�T�IT�� �[�61��H�7�����G�z}�N��#�������]�♡�����@>�W )�I'�����mB�� �̟Q�t�����ȎL���uBp��J��0���+���։Ir��d����ޒ���	fJ��B�l�w������<��bƵ[�"�~i(E�c���f׸�&��彩�o�\k�f6,��m�������KXR��7#S�V��S5������&!����FTB�D���߄�K~e�䥚��� #��Q�&XD���ŭa�ߠU)5�fB���9��w�Sf"_�{�n��$w=���,��n1��"	�$3J'�;k�� �\��/�ˈ_�������C&3}���ė�Ny>��胸H=`թ5����V*�������R6���&�p�:G�J��y���Cӹ�tx�,?�̧_�R� �̷A%�m�]�[�_�K3�Z�M;9�`��[BK��Z�\ h�?��nw�Ս?M���������qSN�2>�症&~3�	�Ii��t��
���^}.A�AL��X �| ��L�L��YD�H!��~�]�"0d��nBÖYЄ��@� 9|s!3/��s��p!F&n�k�*�0�f�O����\#�1�)��H�;J�t-sr�_�,�����<��xu5�D��:G�񊓎��<�]�u��W��Y����m9)���:.����e�Z��Q���Y�$��6�oڌ+#�mY�m9�o�:!8\/s����fD�~N��Kf�|g�a��-�%��YC�-�}�}�M��9��]�K�KԩV�U���E��R��,9�ɬ2�%��kK���?L��mh�s��ws���D�6'_�)�ǧV�hbhX��XdбK	Y@���S��m~]��O�#�ߔPCbnt֢)p��*)��4/}_y�&�Dk�z\ot�~VL���5x�V�D���
{;�u���-�l��j:B�Q�R��M���x�ڨ}�y�66[��ίy�U|�hW˟^���������9�%�>H�2N,���K--��Uf����)ٜ}���
2/nk����ϗ4����#�:T�6U?��F
g�զu���w<<��.��G^������;�	0�g����e{�pSX����,���8�\%�{J�l�e�9_ϊ[GB����D^�!�"HL��7W'Gn`.Xi�O5�0���'�0�v�����ĔXz�j�x�j��ƄԶ��;�;�8M�C��`�[�iz�4�5@n��3�$i��O�<Cc�j�4��+�����!�,E[����_��F�aN�+����
m��]WN��A����F3ٙ��.��D��C�.�$d��1�3>Md0����Н�4�*|7��7-�?�9dt���{;'����ᑇ��0'	��Gf�U��Wc+h��$�n?h E�E3�f	Sjw.��$��a}m�J�� h@�g����6t������d�������9G���_�[Tul�c����KK�WX�F�!^�}򏢅�6�/�2���
����>N�[������{z��2K���K\;h�4�7jL�E�C�x.�4Ê�kA �zq��f�\J/JB}\ʜa�@O��,�1�%`扲4�%��F_J�G�Z��z_Z��0{�}�\�]Z�^k9z����an���\�#����c��Qh���A�W�U�+����ag�Ȩ��Dh�9|_
��x�S
��@�����'������ɫ��(���{?7�>�G���i�=����-NJ\�&���vLȪ7��f��5�
L���}�ttw��B�K���V4�������� �0n����e#t��	��u���o�8\$���(�^���ѻ�DbJ8&�Ț�/vN�#l�e�����Tq��j�޲�>�Eښ�F�>/U:}�g�&1���m��g�4�_������²�����3����F�&����齑�௉-�X���9N`��;O��Lk����Xx�[3��ǹ�;��)s����4h�jR_����/��'"lU����2�M�5"�M��.5(]��-]*���mqLE{L���H��cH����A����0�/;ny�c��ZA�[R����S@���8{머�-|0,8$���%�� � �[pww�w
�$@p��C�N��$4s+��~3��̚�X�Zun�{�w������w�2_���R�ܧ.��k�u�%�C�]!�Jku鵷q�O/&��UAT�I&e���t�{�FjX��o�{�U��^�5#͏Ņ�,�6��:�괶�e��%͏��dX�x�?��*���z�ѐB�C�[i���|(�ߢ�>��x�(�F�cvF��y3�cS���'��ED�i<�8�φ��GBy%�L��u��u��22a4����j�C�Jbh��dG�R��!�BDD�	������3��WsRr2Gӻ�ؘ&
�^�>�&������@A�/U��bA��P=���e�u�o�j�n��C�}Waca�|C�Yn��9�\װo�70�ƶ�2��g�jyY�H�E�`�R�*aq�[�Ee��|�dˀ!���>�F� ud�A��@[b]_�m{�e3�'�c��'j��ʦכ��D���E�������=����{]����x;sYV�ᭃj�-v� ̱�o&/	W���TW��������D�WO��j�Լ.DH%��u��1����s���f�ZG�s@W�WQKS�>*��dȕ��F��ɠYz���� �@r׏6��"6˲�&R3|��\����xh�"� ��K�E�k�k�}�Q�'H|�t�W~X@��������z��u��D�<�[��*oA��{�L+�����z�kp�_�gu��c�c]��%߇�D���ҧc#Ӓre��b\*Tu5�6�t�z'�pwp&%�6�R����޽r<�
�˷���
�/�&��/����ʭ��M�qH�\�s7/o:%A����s$JPU*;�����1';;�g�n��[�Q���C����m�%��9O�����P��^<R�a���H\�>Y���Ie�8)���;2*��E�U�'���{��H�[w���a�:���iAW/R�FO��{��鲒76�]>�4�Ś�� H�<�<��-ǝ��1[�9����f�v�@{���B^Y5��ܚό�o�Ն�]�# (d3��������,�qf�F�QH5������K;R��&j����E��r&/ȕۥ�5/9�Z�閃+�������I���e��B�U0D���X0G�h���Lʥ�3��[�/�r�}ѕ�4�j��zp�n	,�js;8���./�	VD��ڳ����5,�@����v�=�+"?�-�0�5������{�
��Z��Ob��ͻ�Ļ6�2�s����[m����i�e	v1�?�'r�qŏQ?��!�-�b��UԪ7 ���}����V(��)��l��û�c�w���3w�Hwd�D=�2���<���$���l~�|����ꝻKY��s��_E5vO [-�뭗�Ԥ�\�����C���/�-
�p��_$s�j{��8���{vy)��L!wEQX�h�|�yAC���R3mWW��Kdd�:�
B����aDO0��!�P(��<�����ͣ������\]Q�����ʈ�8}$���N0޵ٞ��9&�>�����k��۸����bحwd:u�Z��9��/�}�/�=)/
����*}(߱�lF�� *��.؄+�8&�r/�)�-�����֓��z>���0Jc^sc��ҥ��1jߵK�Bְ��],�,���Ӊ�gK�������5z�/y9k�Aܱ|\��"a�R,ӣX�0�����
����xc�>��E��/'A �&���g�*��!ŝ��eˠO�+�b=�1�;�
v�:�>Ȧ/`V�w�����ۂ�q�ct�.f�I���R<�ċ��Gq�jv�[\7f(���wk�<!$n3j�|&�I�ճK�j����/�b�|�:c��P�v7]�W�s%n)9�Yl�7'��������O�҃|��A�=��=?���s `QA������*�.2��KztU����NԄ�J�N$�Y>�Ŵ�1�;�<D�&�^A�8~@�ڊ���T6�W�!����	��)�*ھ�i�����!UWz�W��3�v��t�~e�Z}R)B^�ˈ����j�PΠψ��s��.��#$D������k/�˲����>�V�\JI�I���zo���QZ�*�?/�	��)Ǌx������N�� T�Y���M�/�4�tg����c��	���U��"�z_���(�6�5���;}R�gp�������O=E�نW�-����k�iK���xH���O�g��.ϻ�q3oo&'��w��l�!�}1v5��X�G��feϧE4L��L&���|��2q�:ױ�2�W<���ZM1�I��WR�������/^��=GG|�H� �qS:�(��:%�j�f�A���a#C>�RF_YgI�� �F�1I=w�^~c�wG9���L�PB"��=<����N�T�؛8�k�9�Z���
Dϓ�}p�3���M�c{Z�#�>���Z���z��9$���(�yt��u���mbzH�奨E�]ڽ{缕������\s>r84���k_�~ݕ�i�-�6�]�,�J�|D��[��oK�&����לf���]gZs>��~�N0�|��ɺn#���س+��}��� �C���q�4��?~��,7
eh�~�[ӬN���e69�*v���r@J��'N��p�EGҺd�I�i�v���n���eH��� ^��|AyuY5�h�r��r���#�����]u2@�tTy4h��D:!'{쬋3?�?����L?�dΚ9S&OG�����ع`Z���-,:�����gBc�����ϝ_2�D���ޗ������ٽ��"������^8�W"z�mP�48y4.��1tl�P7sV<q�H=	/U�(����і����0����㲐8m=S�ڵcW^�=��	Y��o�y=�t�%E}Fb��u���ռ�cѬ�+S�E�@��~��sǵ	%�yNx�w�Z��y	kBk:$dg��S�V��ɪ��@-W)���r5���ϵ1��U���-f83 t����Mp��V���o�J��wM���4�>No��f�k�7�pT̄;pO��s�"���z�Oݘe[���|�����d<iɅ�6��G� �}�g�������"��r��!C�@a;�^�(��/Q�g�cj93_��@qQ��$6��'��L�����e|D�g��~��Q������gG\��)���8�R��\}Ȧ��ȧP��Y�K���*[�S�?X�EAH���f��gr���7Z��,Y���A�� :�ȸ}��!Ý>���������f��6��.f7:IհF"�S����`��]/lmywβ���2qj ����ףb'B�v�OI_��W��u��J�Q�8o�@Q�:*�-@앦Bs�N���O��P<�l��fJoe���$�x2 ��={�6)~ �(�w�6���ό^e`XAH�,�
L�Xw�
.=�<{ �~;��$V7�]l���䤞W�E��R�C��i�W���H���V."�d訃]4܀0����!�̸������5�j\���-g��Ĝ���nA��%7��˝�#���ǽ���E89)�lٮ$���/��p��w��m�o����VO{�3}�o�����|� 	w.�c�[~��7(m���*��_�,
Ie�D$\9|N1�vR:�>i*<畹��n#�\\���~�%�� )x�`�����'�O�_��8~�(���_�����ς.�W0xG;DUy��.�{M:㚐/�x����P�q�*�@]�v��Εd�.���{�1+`����tJ��G8�0+H��e*\����g�֗�.�Ի��p����Z1R2Hғ��vR��:}��k�1�h����Uy�j��V���V�!��\j�ĥD�LdN��cJc����̔W���Q�d��s3�Ih*�(۾� ��]�]����%��{�zB��rڇ����?�G��L:��a}7�w#�=z��5O�IO�(��L���h����Q`[
S��N��[����K_E�Dq�b��V�2,D���ێ����	Ǌ��#��$6�QwQ�x�JuPЏ�L��� ���� �[ 7�]�LMx �x�(u��1+�G��k�B#uX��8_m�X��ʜ�������l4����N���siۭc���g>�}=o�;y����_|�5�8C�!��T��O���Z����`0S�&
����A������eP332�$ ���g���'@�'��e����d�|����A�F���?I��:�4L����B��m-:k.�f����m��CC��X��`nlbS&��~��C�6MɇFN<�ðo�#
��%���ק�tG�����:�ct����g'������OҽK�l[����p-��� �N
&xU���_��|b���gn��.�c���J�2<�4����}�bR�M����.?o����k��ҥ v�3�|pU\�L֍�#a�A��vP1���%��~_B�9�Y��;��
X�����!�ǂcS뉓�v��I�3�8P5#�%�`��.��/��Jr����1#.�f�����(�I��c����o��W��i�KYP�u�W[�6n9���H�:�x����Q��VE�X���%i����à�.M���ZE�!��d�mp�E��e`���ʢ����$m���xx�t��������O7��(� 
��g� ��J"z�8\r�\��pQ�������{EQU��t���X1Y�RjҞx���7'E�	"�2}w�c;i=w�=="^��F���c9�U�x�8�*,k_�V�&�u����oS���7���skXk��1OB��#�s��l_N����L�s�ڤ�e6�� [�N���b��m3r��p�zx��V��K���AW��5�` �6\�W� cs�^k{���rT�hٖ8[����=����!
{u��e6z} �;6t&��;w��`K[�	�*x�؂`9���Cv� MM}~)mZ��z,�l��N���-a6�N�Vn�L����ر\�(��×�:��L}��I�jS����z��Ý�+>ifX�<��Ȓ��z��2�4���a���Z?��Q�5�g�T�|sv��}}F禎�Fo_+�C�/`��Mȕ��)T,��X�~�"ݬ&&1�+6��A����ś?C>�����p5M� ��_!H�{N�\����	
N�5`�Qq
����0�ʞ�8�Y���8����| ՛�N�x�����J��m��9O9S�o���[c�R�Ī����!��CM/������v�1���%]_�[���Ⱥ $ܕ���6:�. �=���d��ov F2�#M����0=�qG�KG�Wd?�"4v,�0��mm���!��4��n�2թlP~%
�{젫���K��yW�
޷� ��������|k�@F�G%1�M�������r���?$25�N"���6��E/N��H�a����:�y	��>�nz�[�����f.c��r?;]|��Bc�li���ObI�jc}1��zh 
�	n���0��dɝ��2�,�<�=������W���NV����VFJ�Nǉ�x�|[����ыzq��z���K�e�=o�f_{���@Bf�}ӽ)��*u���Z��W�/���؄���	7Zfx�V�80 �����Ui�Լ<��K�8n\I�.�¦&-b8-����2�vC ��B���D=������$�J�	��EJĐR��"'k��2�~��R��l{�	V��`L�Z�uA�(��}D-NF�Q`?��� 8i����}�� ?���ڹ�+�����w�����2ݢ���1�� <mnCavv��V�r�f�^�$&��5^X@ʺ�3w4uL	 ���9��@���k��ȌI[����I4J�j��Ѓ�N�js�غ�JDgJ�n�o�k��X����v;(B��-s�����:jwY��7ZX;~��2��F�4sU`c!k [���F��X�'ϝ6{��N@n%����(�nXW��G1#����S�V���O1�����ɰd�l.�t$�ʲ��,�O� �{�e��2ʁS�HR�x�ǀ�ӂͫ�[JW��Y�a�:�Ĝ�_�b��E�~=8C���w�3��.�� ��	C!���LG��l������sxj{��	hߊK���MU]]]'��(LM�������}N�R�ϓ�/�&�� Zi����?72�'��
��@�� E���U��K�4>�=+e��w����\�lc\��2��僯'�Ϻ�1%u�L�u����D�?PQ����7\���˷��v5���nC���V�m̦��-(C��&$H�*���K��GwȖ�.�I���Q�ظ�� 4�ቊ�ho��oKt\��7�GN�|_�u�k 2:�f\Rٿ��{>�����
���4�M5��8����{E4`a$�4ʦ �⢿=���(���k㋅��2�S�q��m�u��i�|�����s��t�˫lNM��	���T��\{���k�R86B�t�q?:��Sp�K���e4u�7�bu>�g�\ە��׻�����:2��K�/ڕ�z���7U�L�_���	����>�G�hq`A���������p}ϻ2�,��|���}�ܰ9L^k.M������ӹ),,�I^Gܢ��F|ܵ���+v��+����x#�����w����{������:�'<�y�k�)�����y�F��8@�Fs��B�\�=1�Ş��h0!
�)�͸�i�-��t�'�Ae��V<��wl����`c��QC���ԣ?1�m2�
�{\(�������\.ٴ0>,{x�њ'�̾�j�g ���:|��"�N��ð���f���yg�-�Ae��[n��K�	����'[+$� "��p���"�3��S�8{���ݐ!��)���. !ʥ��˼�=��x�J�=<4��7���?�(p@�/�w��n~���_��/ώ�؊Y���h\�p7���Æ���Re���1�;�?@���%0�[���F���g�N�q篅(2:��T@ �+ﳊ���#��px�>xe���b6%�8�A�t.��2�>��bى�i���,1��g�ssT�?a�/������DO�1 �i��#�3�i&�����'�hH)R�����q�M�EI�M�}A���m"��剛7AB��Z'0Y�4~�Ջ���y:��ԍ��)�=�hY;��
�>sVazs�,�s����q�iW�*U�]�qVp��.u�~»�=��3@�ͺQ��[�	�*f:��l[�d	+`V���͊i�����{3?%�*�18���B�ЅwSo��[9�x�R>t�{�VgG���b�Pr�D���L�/m�<w�R���}�E�,�Z#�j'��TxGT#��+_�.�(��jZ����mwv+n�ъ��-�mm���8�]����Zo�0�Sަ�B][���үn��F�D�W�$�7���T�.�������X��p&��a�/� �u�p��ډ����He�=���qkE=��t�xv(��F�����O�	���������W��T4sW!rG���|�ߑ�~B�
��W~q{+:�̸E��ha4��Y�����K���� i@BHJ���b=���n���E{��Cs��M��8����k]Z733��ׅ�F�d���tZ&p�$�6���4�i?+�'�d��^���e�Ī�[�ͪ�ϟ���τ����_�퇨�Dw�R�:�l�g�Kޞ�?"�A��Q\�TtT꒕~�W2��ʏ��O�r��pd�F�� �e����0��c�����D'0-��YF.��/������: ��`H���������T�ކp���&�S_sgQ�ͨ]C�"f�sj|}L�䠫Ca�^�Z@�p��[��Y��=�M*&޸uʄ�|:��zj3�}�+:���/8޹�|�h���!(E�a^��c)W��k�{��:у����e ��u0o��3"����a�J8�yN`"�e9�lƫ��ص���Y�d�4���<�w=�%Uf�M�='��#!k�\�b�ʷ[��0<F��_I�.�t2�N ?���uW
��s�d�;�S�-=j�O����]���?軗�X��,�H��V�e0�D�����w��V�Y=|<���y�pжw� ��/Sj���l�<��n�� 5qe��֦��}��f�B��a��j�D,4#��5	����Ӹ����4!�W�,����K�_�'=R۫��)&ِ���U��	��*�hU�Z��C�A.y]���b�������_�
��,.+KNI!����
{(�{rx��o��mm$N,-��\%^\�Y��$�fday�O)�Km����%�o�CT�ug4��}c����~"\���	횋普���fͨ���!�~�F�c�������k���b�J��wg�\����o�4!Tj�n�?�>�KE��ٸk-F���׏Z�N`ز���&Wܿ�Q�5cϹ;�p>9ֿa�/�!����k sEV�)Bz�3((�\:IpGVH�:3<#Pf�m�m-�:iQ���h�:3���U����u!�p���yb$^��w���v�t(0[�aJ\Rr8􀴞}iP��u�J��ցaF�po����0����dk��
�V��x�p?����"�T�k�:ղҭj�s���Y��Ž�Lu]����F�4������ִ�Lq @m��pӶJ+���S�lNj_�]�v�sP3����`��ىA]ջ�Ʈ���sԷbA^�ݪHї}����o/�H����Ԑ����� W�u��z`� #(dwG'M6�2�T]
*ȁ��f%z���i��R��ׅε7޼�y�h��Z�����ݫor|�)ӓ��$�߅���1��R1Ǟ=�n2+�z�Ђ|���/��Uբ�/�gM� �Y@�� ?x���2<<\m܇=���N*�$���O�$vW+|>��}��w�y}[]�9�8T�ɼc�'��J�psa;�N�e�.��8ve!���(��xQN���������ώ6P,6aY����'�sB�y��lSř܀�r���r�2�K%=��N�Q�Z+S%D�ͻ�d�f8{����m�k�֏�����HV�X����ڕ����X�����(��i%�q��m|�0Z��N8��+/57�����n��L�3g�-׉�4s�2D���܉b���yJp�t�s?I�/�2�kX{  Of��]A@1�G�b�E8Y��q�zӝ>�0����/��[��[�&6aYZ@�Ƒ0��se�浭	|О%��?��p��[I����x�Nz8)����wbBv{��@.��U�k\�E�W�<��l���
��g��bJ��%�H�Vy*�L g�t���̼��}��(�mB���؊/\9������^��Vm*�{L$�۬H`����f�e��Ý)��Q*%6�A����K TA�&�.��>p!���~�n4Xa�=�+g�ბ��=@��KS�ə�pss���dB��[Z����@���f��X����j�K;K[���G!�***T���f�QR�R\��ccq��EYB�_�J�)(C�8Y��Su���"R����H��p��y��������n�GX�&�'����t*CL(-�z
�~rx�t�"���T�x�A2�	I誻G�+�G�U����MK1�FN�7Q�G2�ڊ�Eԉ��� L�'f��|�ۛ�R�U�O�tJM�G�m�Ƶ��>�C��N�`}����Q#(��H���.��(���7�J���Jk�ɝ>(o�F�2O1�TҊg>��m:u4���nV1kX@�͕ݠK-(�g�SfF>k=��qm{ꤼܺۺ�YS�v��_[��-��x~��{ɕ��c��G�q�����p����4� ߮~d��T�y����"�
�q,�L7տ����h`o�m?_��+tX�����"Z�cӘ��V���>��oD+t���W��=�qs��e�"��V��Ƒ�7��L��_��� \����5	s�nj=����y䰧�4?�?q�M��2*C����R�$�u\�(|L���X�\a�
a:���:}0���16fq�H�7�f��edc57���f���677o��{*��z��M���imޗ�GЂ�&-++���Z5��T|����JA4p#ǥ���Y����U!�Q=f�~.��v��Ȼ:�7h��߭�,~l�߿�Iq�7�*".l�G�EOŲ���ѡB���Y������%KjdG^�r�C?�4���N�J	7�|	)bnVx1�à7)�Q��g�咢E郜��،�ɂgTS�X�i�i�������A�3�{��P`�F:lV`��	
�o���u��1��p�B��3s���^ ?��:4����[���=0��?�/�����D��R�P�t�Et�9`Ҡ$%�D��E����J��<Z1m s�˃��Lxt���e�e��[~�L�Jg�0�-}D��2���V����Fa��+��J]���GV�ָ�<&���!|SS���x"Ʌ�\���k�; `#�x��4���̫E�Ǿ1`Y�|�C �c�NY��xM�I��]�����H��7Q;���|5��28n[��`?�˨�R�7Yrn���EU*���X���e�H��u��!�-���Z�3`�$���KJ8�/2����9@~l�m��y�e
{N,.�p�J
�*��̕��q,��BHX�9�\�
�BM6�|��Ś�U���is?i��|�ҥ�NF4$tzv���Q�+�4�t&]jam��+'CW^�=9SF���j6%����rBz���f�3	Fj%��� �syl�,�(��9���`�J�f�n:<7Rtu�a�p��,ln�C�~�n
< Z��#�$L�g�5+< ^��7 d�w�qqC~�:�9K����"���]���Wf��wh�]�Њ�74���ػ�R�������s�&�S5�`��vsg����t�zm-]_�k�/�����sړ1��7I�tG�zّ2E���~`�k�]�肄2�^�SF��̄�S��3v3ZhQ�1�����CÍIt�^����K�$�(����� '�DB%eH}�Z@AJ��<M�~-�˦6�����S��<0υC�r>|��=��la�
���5_hܶ:���ay��l<g�[Z��nZj�X��u�3?��(��q�53�EB�`l�R���B�4T.)--(.~� ��|hC*@E��W���*r�s��������'��>)�^����R6�ƍ�2#���A�#""�_�?�(3�|���,k%ϴ)�N�sA��"�M��Ku��e_5[>'�fЕv�vOΩ���,a%k~s�Fﵒ�w.k�f;�\W���&Y�u��s[�p��
'I��X @Lkn��`N���p�|�y_Eq+qsY����GK�����=�^lNӉ<L�&�7m�9cc����2e��r����hK"���;<���Z]�U���I�v��
>�Ó��_��3����fT���L��"@Ycу^�Qp'(ma�̗Xҫ�����U���EZ�UIa�ikl�]��9����Us�(��aRy��<��$�R�@c��4�9&�H�k����  ��QW�6��ɣoF��ee�y�}Et����yފ���w���dq2��X��6�Th�o��y床_C�kؾ��OCxp0?�=`�����2<�ZmpЭI<�����|v�)��o���g��T�e�d���>��uV}���xl@���Zv�y�ͳ4����0����f���>vXAy�"7�����j��aU�fqQ6g�I�����1��6`\\r����)))ң�Z���GK-���x�H����a�|[�p�8mn��0�G�j*�>G��g���ztW��5���G��?�a �X��8�`��ƛ��Bߤ8�j����:<{���f�v�9oc�ڝɁ��pB�{��^C�L�:�a���!4}x�x�2���;�t3|9ܩ��1�t��0�k��nk����Q8���ͷ�H�T%���3�.<�)����}�Dh��-�8�xI�g��'�%��k㋄�����F/4y� >0�r���J�t!	,���q�A���e��YY	�ج���8�+~��e(�����;a�!.3���1�7|����/)��B�1�c���˙�`C�)�cs�Tq�y��z)��6�;����uʸ�4*m��eI6�q��}.7ߤ���:�p'�ܫ��)+�KI6n9#��BpUJo��G[�0oדwDv��l8���y�䄖�$�벡�J�0꼇A13���NV�3�Z�W'O�;���S�9����������'�D4�)9�	&����?Kp�
â��6��	�Pg��_m����ׯ��)�<�<]��KM8���*Gc���zEL(���6=�D�µs��]�|�Jv7:��_[7bT��J�̓����o�!j�VG��ig��\0-*6$��(���{���o��2�Ww�!pw$6a�4bns����h�D?�$��X֗E�,=���-*�:�`�'ͬ�a���J;�D	��w��p��y"�3=�	�B:�Y�K��ܮ筺�@{ɔݠ���޸�~��ޥ�y�l���y�ԟua B*z:�V�B�v��s#o,���I4��11J���ά�O4=�X֤�a�'٬d�43��8"��Ѩ�8�^`�o��	/��z3OML����<��r�0L�1�4��_{������<s��
���]w7�c�����f+������/é�?w�쨃�Ш�D�%�����m5��Ai~�~�Y��6�����N~��66e9^Ĕ��Y �o��g*h{3H���[i�	muzo&���Lb<q
�@�X=�����Ԗ�7<��"(�!�E$F���><<<���x��9�夨)�Iplj{~�Z�3\Z-�q���)rg{r�J*�~���l~�͗��Z���f�&I4�h�ۉ��������g_������9�6:�b��M��I��%w$|��
��|"ƌ"֫�q7�3I�
֖�)dRB�m�L���Y;�<����	�墔H��Դ������Oĳ�ێZ�ߨBv[&L�n�����݃NJ�K6w�?��l��m��mی��zX�*6������1���N�~��y���떼��X�+��F�sJ.{�E��܄��^mQ�H���"~�W;�6��.Y�s')����V����c�)ȿ]:-�Ïb��6�>�`1f�?�W����`"�rF�`��M�z�LB�����ϳi�ZAC�~u��g0�@6M&������RE��]+E���XCk�]J'R⚽7�K��*��zX6^�1 <�m������d��7�����"���f~�O.=�!���WK�{�*Lz�-�ƳXD%ϵ��Ϟ�[����b���78��}�\�YX����lc!4z�Ŀ��z'BaF�ns��'&[���X}�Ƨ���q��pq!!��]�w����>�yHB�����oUF�i�OG�?�~*J�#Z񤠣�;��N�	� x��w���B9*�RAQq��;22���V�K�Ա����W��Tz�Z��)������kff��˗=%}��(kǳ�w�BF�yX��3Vq+����N����wː����%bQY㯵�q�x4yЧ��$̀:��L��A�F2��ª�fv��7M�����_6���>+"'Z��_5(���ቑg\""w�ڗ{Κ��H~�a~r�/�P^�(�]�e�	�S[.���Ӽ�l���ƫ�E{�+�b줊�n)4
e�@�ݤ=>I�T�ʸ���ި改2U7�`ϳ�"c�~�ȳ<zOܰ�a;t�,/QG�$��f LH�~�S��i�Ĥ�2�;�������Z�NM�		����A�`���=V�%��c��9���"|��B�&p�9΋��
�h;�9�W�SxK�+�O��IN����_�NŦ{�O�!���^Q]�ǲ}[������Zc)���ؑ�����^��}�.cn~3��xs��=�Ƀ�R�8���*G�e�H�^��$��H��a��It,!B6���W��-B��|p�; �����I+��"�v��L�/�;T54q\H��s��(c؜'�''��%��B�y_�NT$Kp���prq��Y|�ln�+()�sh�dW��N!"��:k,��|m����D���4�;��nu�����l���_썀,Db��L'��w����u5V��17"�Nk@�$��C������+9��T�����C����AL���cjw ����1J�Ef����~�_x{=ݞb xf���a��C7L��t��:nT�t1��o�4�-u��NE�β�ϖ��T��
eDblX��I
*F������h%���sG�snb)3ssS3��?��FA���7��٪��O�6G��[�8�a�w������<~!O=���
xu�������(��N��u�}6[�Y�V^L���k�\��h�?>���Pr<������a�x9�ߛa������e;���Ӏ��F�^��;��Qy�y�*
��@@����.��Z|�/�S���|����*���XR3o�n�$-=eY�'m���Dtߑ�r9���C�ڐP�?�H��F��߇@�ۼA9׋Σ�tt2�@�HQ�x99δ����i��ᏸtͼ��o%�)���.��md�Ç��2uG\�X���u(� P����Y��H�?}���K��<�b6^j���=�U��/Z���I6���v�6]�X�P]x-��l�j�1�ԫ+OXJqjh(���=!�Q�dum-͸�����	�hŧef&��["�#z�*k0Zf��:�� �w?ȁ�h��M"���ˡ1����]��?i�fo����m�n.u3���ƃw���<�ξ�5�<�f�����q
t�vv#�aU^��(UU�{���7w�+�X�'t�)9����rh�"��g �}���4�T��~�v��B���
�Y��j�i�ǯ�����;F9	�X����&���7�����C�hqQ�E}�Jㅄ��c�,F��~6xҙ��w?2�WM]=n �����>ǲ����\�0��IKK�%����5y�I芌��3a���Mh�<���q���䁎���>N�v�ebXYZ'��1�f����dz�.[��[.��~ͻY�P/��/���Oϫ.�_?Ԩ2�<X�w|%s�{�f� ������d�����T��xLoۛ���<L
:|��ݷDN�Ƈ�ܝ�# �S���zuM���� ��l��vG���r6����7� ��=絲�4 -��K-�:}�w��	�wj-�EJ���J��}��Bki~�xH�O�ž�Ԉ�� �ܼ���X����U`,��D�1�)�a��_� �P�o?�U�.�)�ȘN[d�!E2l[5ă���� �M���pr�̔��H�o3����[vB��5V�{۟�C.���0��2qq�Y������z��q
��A�
?�r�"�剗uJK���xa��a���j�:�3��z�	`H"��s�r@��~ǫ|��=*D�=�^yJ���o�	����Py�Fb�+�_;{v}:�#[�ɰ* FZdrp�S[��#�Rllx\K�W�D�1�%V!s7������/Q��3��F3���4��+�bn7���(�L}�@V)N�n�'�Jr�4��x`����i���}?U� ���
Rx��}��~�w?A��;X�O�@�$������F�?8��U+)��#H��l�]�mϑ|���?�C�MqzwՕ���3�b?��.H�tq��ovϏ�[/�Bh	tg����!g�܃�Cd������y{q�����Q��kx̜o����R�I
#�����?÷x�b��kQΟ�M|4��u�Y5�ʱǴ�N)�k���o�tS���&���"�H>j��u����[�C��*�d� ��T���O	Eť����x~2D8��m�N���4���!B�nY�s�{\��9)��i�gЍ�c���L�!������S=���w�!�r�nbK^/���J�ўaS�,��/���Y�ew����������pDVz�d5��� 	���1�6Ы�,绰7�D�Ĵ�s�4��-�>w����+/�Y�7K�/���
3!������� J��o�&��M��íi�ɔ�˰��W�6^�}0������/�r�w�&/ӓ]�S���.�u�=��vG��yǎ�G��xS��)��vsN�$��K�_�'�􈷭~�n�1�;a�˝�V���B�z�r�]s����Vu�&&&e�b�� �+��+���+�486_ r��~� �7p1�;��������sj��=X��
�iv����j���A�XU4��[��jg����M���ѧ�% �~
3į�
�M}!��C��|5���1�r��c�T"���\$Ҵ��zbB���Q�8�������7e��`����W���=o�.t9�i9�o��1�E��5�Nn�$��e#��9�V���"�����u���U�9�.���B��n#��%Z8q�����?)N���r��b"����Oe���|�1���v|�ŘwѶ7�Nb����i����%��6�j�v\��}U7����=����b�^����ؤ�s����"�1P�G��E��q��',.@T�'_�ݽ=��8G7Yp:�8V�;��s�Җ�.Y~�N�X�h�-��j_t�ǌh��8����?�9%��	��_m�~�&�$�8j�	U@E�Eԙ�ౝ�"��rY�H���}� ��eL^,�W�tq��P ##͌)<#<E�٤;x)�1:ն�W��o\Ԕ ��������%W�'d�Z3�w��ݗGw�U��|/M���);��"�;���V:���MK��`��Ϭ�<#�F���$*ب��^R�G��wI�ʅH簑aLR+j��v�~��|�W�G��s���^�r��k��+�߮�\��E�Ѡ�כ����t��#[�w
rY%�1`��r����oV���.b�D�o(�w���[L�6����٥#��,:p���Rd�M��e�kS�2}�Ŀu֫
�l
<n{-<S��0�A4֘��
D�y�Fš����@�ꗫ��wK'6�������Zv���f�9h$�K����Y�E�v{[P@JR��n�U����!�n	i�Ρ�[��r��!���}�~}�vߣ�qz33^׊�ֺ�i��7�KE��F��IG���p��E;�k+'ؚIA �1���=\��y� ���I_Ex���K�NW�ye���:P���w#	��u��嬓�fNx2~����8�,���3a>��U���y�|e�S` &�yN�[��r������}.�W���.s��*����#�/�Tm�?G#���ԗ���@?�%�{�ZP�~���p�>7���X�"-���7sN��r�'���+�<�^��>�dVl�fx����o�_�z֜z��Z���|��2�X5EDKE�I��	��o���+�,�,����˚��b���LN�HC��*dlݠ���E�D*�-
��L5�]�B�nAo��n�T~||Z~3%�J�R��7�l˗6�2� U>��Ð�r�
G��3��4�rR/yL�Gaوa��Kʂ]t��_�<Z̏	O�1�J��Ay�D B��pOA���$����κ�$'���ş��TQK�e�~��K��������ӗU���HY��v�J�$GS(h|hyש���@=�'^@]�F��ڳ?XLa�VґS�I�*��g��'������=<y��F�WS�*b��m	��x&^��U�:y6�#�+����ur//-�G�߮��/0˙1�{y��$�����Z�����A8� �H��Ar^����*�M �%(�S�k˭����I�a	�����������c}���G���ݪiw�V���	�
��K�Ǌ��}��=<=zz��KK�B��O��3���U�U;�K����v+�	��t}�H��v*"u�i�a^@��Y~�G1T0c5��R�w�M����7\
J�.;(Dw���4�EбJUr_��A���eB �ޙ^�K)I!m��3q�7��A8�u����Dux�)��÷W��C8D�rq\�9��rq{�����4\� �� �h猢G��7lJ�\�O�������ʤT�(�C�y2�@mj��� ��n/?W_-#����@��8��CGYq�w�o&�iy�?ۂ����y���r�n��\O�
sN�Rݯ:f:$Ș�a(��x��`�����ҶK�G�
��ly�����y5
�ܑ�4oJ!��^�K��e�,�{.?�8�`X���,�f��lV�W�K���u��;߻8��UP�g�LU������̡z��ʺt�	f�����m����⠐��FQQ�n�b�e;��Xn���h��|���u(�n�+��ow����g۷����EF����/?�:gz��U��._�p_e��������)4l�-��'��F�kry�a�U|��ϛ���M:�A���铉�[��e��c"���Ҧ3md�F���J�(p�@6�.�O?���~ϲӰ�Ji��.F'q�B�h��{^�2R��jz��ZSҼu�_���a�0��jh�P*�Fڰ�!�_ÇF����ݑ"6r�A�d��]<�H~ �kH�'�#�uz���N���L�̣�	�i�Ί�ڱ�@t[i��Q�	�۴��V�7�	:svc/�I~�zJi�9i��l��x,c�m=LH<�W�#j���(cա�) #�2CT�f�f�IY)s�2%�B���,�5ε8}�n����
A�������k����ݯC�&�~7W(��k�k��Mā���f���v-O��Aȁy����0�R_��<���J�+���<޵<;I?ߛ�����9j��_k��/b�"$5������-ʿ�晛�������^���1J�����B|�<�\���U��D��S<�hc0�����U{ά\yx1�	~�-��,gv�&���N�A�4�|Q"	)��\Hp�.�#�E�����6�zXF-׍
��\C<�^yŹ���G���@G��&���T]�����a�Q���KH�y08�_�~|6��3���iWߗj[�6`(�U�̗t�|�t�,Tܲ���E<���z���)!���O�f��z�B��ɉ���>KOj��׵ܐv/�0^��Eg�<�"te��:��ҭ�̔�Y�p=Y)���وdŕ�,�qƥ�:�nM��o�a۸8;��>�]Up���D1�h��́^Z
��-a�az�l#{��/5�I�ʇ)M ~������J��B�4@��J���%>>ALf�	|M?u��o�f�%5�D�<ȑ�����/���ʭާ>�;y�?OY����<���%���>�������:�1�^��w|f�)���<��O�?;�����WѼ��-G4lx]k��]U^⊅��o����,���U�����q#��wݪ��x�@k��EZ@��uM��q�/_WFj^&�i�M�^��*�23���&q���&E�bY}ԼBb�lX��M�T��+d>e�+�&t���֢O�g�������zm�f�~HuJ});i�:���r�Q�߉y�k�r
�ρܧM"�$���������$��|�|�>������`�ɒ
�W\���E�#��E�������3)�����u7z��F�S!{�j��c|�6Wj�QgJg��p���$��y��d�h����Cf��p�E���~�Ps�3��8@�E�sKDk�<8?{�73+�X �����roߢ�=t����V�(����V�~�.\4�x$>w:���[p����s�Lo���|�J�
R��"��{mu�s�ў��^���������.�xtv�m����w�ữp�p@������j�{76q�s��(���hQ�:�'���kAhC�.�⌦�?�Z���N�e�5*��{��s�X��5[��<��x�$�<��VUOM(�/�m'`j|M����;�V��\X�39�ᠬ����<�O���'���U�}�*�j�6�x�u
5�so��,W?bW��}��_��N�y����L���t�����=U�,3�̕�,ᖎ���[�P�~����1������b��˭���'�x����fٙ�:�n�jl�NQ���mmf�@�ݼ�m�2=�!�!4��IڨYLM:��c|�a�AK�+(\����4xH�[�>��|������"����Y�Ɖ}(��u�aQtp��bE�-hty���neYG\��UlI��R}{>9t�6���rj^���;��u�i�>2�ְJ'P��ʠCI���(_:��Ex�����C" lv�w��բj��i���dsz�z4w�N���ͥ�R -��DIr7��ˁ��
��'�����w�+ ����N�����&����_}����g��-xɜ��,����#��bȸa�\֒�H��S���7\�A�o*�����4O����s�;���)�>I�X�?D{4��1�\�XoDC�Nr�n=2Z��� ���d���:s,*��B�h�ݗ�� w*�9u�%�i�9���9��EyeKtg9�����CT�\�Vw����04�ѿ+��]��õ�CJ�L�U���DԒ��@Naؠ�a�a'���#�Y/d��u+Y� jPp������~�}%36�u�UL�
bZ�s"4��,,*KT�i:��|��<8��)�/_��Tph�,
��_*�?V�a�t��g�`������r?<u�ˆ�����U2{Y��<��?~E��Yg�����q��o�$9����U�]fXz��I��k�c��_>�e��L�wyWG<i��(��8�m�<>̻�%��M�������t��Z�Y���l��*���uA�b;�^�9�
��W%pk�N_���c�o�o���u�Lf����YI��|+�$�o4	]�^Y���풇�0���L�P��<��F��~K&�)��Y`�}��V����'�E*qrٚO��P��&�S��T�s�[��V�~����u��s�
_'�$1$b��/�P��y�\�y�7
s�5�b(7��M���G�� ,�Y�i�����I�ɶ��8j���˹����w�up��68�W��܏#������I��h0Z�s�['�|8������O?׃���cp2X9 Y��uv��rOh���½)(��./�/���"��_�T�Jd�"ɧ���A�)½�I>i���Yi�5�8U���$�c��(��.�ɷ(GڽO�'�<��gތ7A��WB-�P�H,��v��.%K\p��82b��W,������W0����ѱ&�%�4�k�X�`�I�X�J��y��%:�M�wY���ڐ2�l�PjI�`�ףb4޲�yetBs�w�/�u~+lG|Bu|37�Qp�,��PQ{�(Ț��l��078�-�����~�XX�j�ޥsYRf=�'�qU�V�������ϴyM��B��i�~��TF捒�;n���i�#~��t�~�;�G�zQZ֏v�8��L��%����׾[T�}g�T��"M�6Z�Xױc���ce�	�?mg�P/\�wo��F��gE�,
������\�
�O�sb����+�%��dk�
Ҿ{+̡XC�u�}�r	K�TX�9r��f���C���`���+$)��KO�m����!4������I�+������'7�Gi����t��)1L;	R�0��$3�bJZ�)�T�ݿ�P"c���os�]�1�k;9�5����������-]��
�k�����4R�F�f���.e=ē�qo���n��T!!*:�7M�/p�1ԝ�z6��H/����2��"K��6c�r(t�T��Vy�M����D�I���X�Xjϫy�pM�Y�k��C�:i�w*��Qmk�d=�����)�}��,�ï��d�a�8�/�oA�wِ�F|����h$����w���s�^L���݋���	-��,����Ͳ�	$&`������gBC��8��p�C�Դ��u:)�ˆ�x�z�^�O7���?���(f���Q�3J�j݄�?q���2�nlS����^���L: �Z�$Q�wG瘐0_S|�a��5S��^�_�J���ТM����cRR�-��7�864y�#u�����̤�>�,Oa2�����M����o�~&����w��A��	�(��휾݆�kx,�Q��#r����H��"�
wF�j�U���0o�����_C�	[�׮wCJT7�ȧ,��;��>����/e�5�K!q�Aԑ�}g�T�����jD1�
��p>��z|����8��R��Ms	��xVJ�9<���� o=��ەg��wɇ��_kZK�]��4��\ճ;,R;� �E�Ϩ�XW�)O�g��E��<q)Q��I�v�x���&��MTIH@@/$������ק`aQ���aw�u�(}�`X� �E�id�??�P�9�R�OI�
b�$��rgE$dVS��[N��Q�:�?to$�Չ;��R�P��9z�)mV���B�{���S|����z��#Ju�w��fhf�Nj�wޗ�r�5Zq�y���R��oo$k�����s
�Ev�f�.T+�n��~���}���f�r��ʒ�����ih)D�P�J�>ۆ�ޜ���� �R|�<��d�:,���}u�T&�[�&�,ν>s&��:�Hf/-Ʞ?�t���96A.p; i	S񭨬�IM-	{����.�BGG��u"w��ڮ2O%l�H�홧����t5O�J��)

�5��!��5[�Υ%��Cywߊ^��nƽ�r��D��5V�߾T%�O(�v����[�1̞�5�W}.���pQ�֑x�J�K�/TGk�O�k�臭4bx���A���te���>�.��xȤ�Wlsö��&k�[���D]��sK��Ս�52
����*١��[�wڲ�7J��A��,r
�ϟC�����j{hsDR__3�(T^����߿?���:!&����E���<c�?xΙ?��E �KV��v--c^I��{����m��EK]��f����#��0�֡OG�q��&(���t �R�@0]:��N��x	V��r���\H��������	�g�h��&�TϘ;�d�����w���o��������Ǣ6�\XK%U)�Ez�b��Cw�Q&t�%<�OӞ,y¿d{�?�^�||��%&�0��j�Ӛ�J�2�D�g��p2�FICӍ�ź̜�����#���Aʛ��j�`Kąd
o��I���,	�����2P�^l��9�˾1��i�8&�5�P��2t��q+���.U�_u4.��.U��P���s^Y�$�9��u8�\'�q͆#��N��/���]G�Ҥ�����3S)�3�nHM�c8X�'K�=}.zB=0�Y���|m4�%y�G��T���D�j�����z\i�������⃞�<��"�?�ōI��\67�cBzb� �������(3i����[�2����.㊏O�xmj�9x����y`��A�N]W���[���QA&��z���'&�����T	2{�����l2�t�*)��-��+�+�a����V���lߐ,���Tz�Ą+j�!�/g4d����4ʷsz��j��*�|�.�f�y�l�	SL�
�B�܄����N��]�`�~Y2E���U51Ʌ��"E''3��z�R�͛7^���7�>�Dނ�Ed?-83N]�>��x���TQ��`[�PWX�0���a��c��fs�4��XTZ��]c�قOc�q*)3����������В��kZ�nЁf��R�#Gԇ��!�-���ND{�����L����'JpO��@���G��W�H�(^&�6��V�T�m)���m�s#����㓕[
���0��K�ԙbP-/���4Z����N���e�R�#�P�4�oO��}qБ� %����}�9X�m$�V\IlllE#�����:��ML,�N���#q���z��2+��;�o�ξ}�\��x�$-���J��ч��OOW�d��0�/�V�_��5�nX'o����x�R'/��h�Vl3�q��}�\��A�f,�w�3�*�A	�R��Jv�r��̐�y���a6��dX�{{�oݎ)�5Nav�;8�(����`횣�v�"�e1���,���b]fe��^7�"T��oi+K62I7��6~��R�e�T�{x��ƶ�brkN+�����Y=�]�W�ҹ
?n[��86���Q�IqR�Ά�͘Na�G�gUfcO8�gX�՝��5�8Mn��P7W+�;n�P��Dj���Vk�c�`���!��"˷>��v�J?o⅐�t�Y�9�|q��˘9qH���\�޸Y���������U�R�@`��X�k]W��ԩ}xt�ϵ��U|��hE�Y(�'16}ҥ��n`��C#��v��rP �Q�򼵬�U��������;��f��Xb!���Y�!�F�q����n�m��0�ʍ7HKrU��f4_�2ăh��Daxm<��M��3����Խ�XP4�3��D�������-��R������ˆ��kΝ@u� ����qғ_lr{�&����4a ka�P��<�����-(|�n �Jl��#h[�ZJ�,u�f���a0������YEU|,��|O��;��r(�=�M���
�.�"�Q]��#K�G�I�s�{�<�����ݡ���`K��r	��٨,^3�_z��3���2��A(7��T�(�>sWy�3��~ 7���R��\'�u���ެHu���ֻf�%�q����m>��J�#���Y�����3����C��D� �ƭ5��;lB$��f�&LԌ&���U��ކ�/.77;�;��Sb�5`y�Te�[M�FsÚz�u��RI�m���X%su_ȝ�������+:l��ߐ�:���Kq>�Q��+��&O���As��g�ª!���F�T�Z��+�ïJ`�$�LQo_�6mA�$z���f	�m�쥣Wb;��׭�XoΞz�?��k�t����7
�ܭ_�<�U���6���w�����%6�$�b��˶7\Ն��;'uo�;I�����uhV.�ϒ��<)�Jjh$*(*�#:i��v尞�fAiA�?_��[4������ q���17������o�S��l�G_v�8h�`���Fj,*,	I����F�+~B>ɉ�u���uУo��U#��Q�X�e����X��JK�&%A�2ē�_�����=��F�Z>��gB��9.'hMvK*����l�r�ߩ��
NQL�;�	#	��MJ��[=�j�����vg���O�wjZ.T���^��S�⫛\&C��� I�I�V�0�4��C�Q�d{�=�{�]b�2����Ԡݱ$ŵXeO�x�V��0g��or���q�������������!�w%l"l/�"��ގ.�҄r�/�1�xgt�Z�-�	bn)�*��:������y$�L'�gM��C��BW�W7���f�ʙ"��/_��ML� h��ed��)*)]5@��sZ�^�}{�m�>"���y{�������?)�VTG��ѵ(��=>��[���G����T~��.d7��ܟ�����f욬�ixU�I�覊��ФL����aP�2���"��۔B��2Nv���M�M���p��;=c�5�7�-��"��H7�?��ڷ;�"Uy�dѰ�k�ęm��>��m������������*F��HA?\{Ӫ�z��`P��Qu�c��%����o�l=��iؾ>}��+q��������`�ҴT�Ӛ �W*��I��ʻ�\r�ֲP)b�u�HvǋӶ�f��՗�nWo�=��LDn.�!�*���5��2vt����Ў
�Ж��N��Pb[b
���mץ���������rB��� �F�Z�U�u��4��>=H����2�}����':�{�SE���qf�8���Cu��y-��^f����D�VVTx8�1�!���)������L�<8���B�fKj�0f���Bź.yh���� �r6f|����z�S�Ya,%Yٗ\بi�w~�o��~_���CȷU��V5���VS�I�pEu�e����l�P,�x���v��%�0�نW�S��F݌��J��6��:����ǵ�bcaͶ��aF�1�x��D��#�(����mj�\����4E�\��`;��7��٥?4���:�I�.��k�deLK:��j��zі��LI�c|�{QG��1��z���L|7 E�Ҫ�G�t��Ɲ���p~@%��\�rW��DN0 �^Jn&�uJZX��O��ﲼ��c��2�u���0���˼�N��@-��doo�%**s`@*��eY��a�1o3WqP=X��d0�׿���|��~������a���b��Hd�����,p�g�j$� �5%S1`pޘ~������*>i�� [�q��l��q#R~�E�/��
�ʳnTI�q ���Yw�|�W�ZĚ$�=��Ƣ�Rr}X��y_�eh��r;Z��|��"�1C/��m8��(����m	I����rn�a�� mzx�m4Xu��d��f|\�%r�/<	�/���1o�-��y����T�z۫ {|/р����v22=�ѰdS�J3�`?
~�v�,-��RbXZ�ʋ1������.�G�����S:5�S������Z����*��":5B���KJV��ZXX�%:�vؾB�y:�+�$�$�/�x<��m�o����B<xS�=|#��,��e�µ�3�p0��F���82�f�j��:)�
/��o�7�~���J��Klp+��>翀�%%�؝`���2�u������_ӂ(AMbU�����wԌ�	S��<	�-''�9�w׍ޅ"F��v���]Y� z�7�^gP�'*�%���.��1{�gKf[��{���k�%�߫e-�t��w_Qb{�a��XVjZB��,��ʥ�� ��܁.Z�����Q����jw���Q �oD2Mvf2���=n՛9�]�9���}��t���@!��LnffF�HJB"��O/*:���)==�$��P)Q8�\����ϞYX.̝����qzr���O��v*���%殬e7Fغ���)Z�X$oӳ,�~���n��v覧e��A@vs� �))�4:Xu�����Y��3�` �r�l���� 9��_g�e�H�3�����OD�4�+y%n��k3ǎ�{r	���E �SH~�:���F��#+�MD�d4���c�m�(��+��G`|�}?�["�ˤ8K���w�����%GQx�3DN�9�/z�c=�^�a;f��'����ri�D�LoUBN�J�q���r[^Mo��H���|�t'��O��gQ��&{�G�>�L���ͫVQ�r򭱞��⪩a����k8����Z�q/���2�Ȁ�����Dvܹ���lZ�U{���4Y2Α0,�{����~eC`5�����d`.��c���jm36����<��+:��-���X4�OS�N��U���K��=�w�<{es��홢99�7F��}����-P�b {'�Ts7��ęrhmbϩp��T]��!6�E7	8ވ�o�sT��(��H=�}C�e3E&����7��8Po1d�+ޝp/Ys}!3��������ڷ�5���t�:?���G�b���r��:��B,��,E��%-��|z��l=1h7,�Ý0�"l��E�����r����Y �`#��t/���@^��x֯����Ȳ�$Q9��T��Yx�H��� �A��v�/��Vm����v���}���wn�È��%O�q�V� ԟ�P}�Ъl�uLJC���,�A�(�D`{���L��aW���0j�^�1��`�~˷����P^�zN|�r��7�e4���:�d�0���u%����9����/�޻'s��nI�� Z��m���*:i]��%�9co]�p��P�m^J�0"�1j��oH`I��>�҉�XQ^y��7�|�~{�iqd
=.����AJ���Ze��fs@�6�6����f?�{��u��ƌ�p�}�pu�q��Z�12nad�k�Wm6��	�|F۵#���y[+�=�=.Ί㨾��L?ݩT����J(Ŕâ����}-���zĽ|�|X���������{��D��4���{iZ��R��˃�A����	�R���އos�����ɯ�Z9�XE`��!���K��:n��)�,��f�۫�C�2P�Ҽt_Y�]ݵ�0VC��4x^��=��^+GD�:2w���6E7@C����7��ǒ߃�,W����E���8�iEqYe393 F�������������*�=�2Y����Q�\�6[li~F���>=���oOf�A��.{݇~@�-�@+�V+t'�/>��a,���?T��	5$�Xƌ�V����%V�M��]��K��'�AA��L[�k�k8h_����x�[x:Lq'6����������ZX�R����G�d7#a��!���8��p�������9l�����R�֤�ڥ��l���uR�C��8�����2m-T����E��@q�������=]%������3yLY�(�Nyj𜹵���PrE�"�xx�c#w�J_>��9�ZR�N������8��ԙ�E���#l�0{5;/e��T�*Eʹ�K=6--��k�Z,�m�x�j]��V��s��Kgz�7oې���t4O�[#.
���e#'�X|*ʕ��D������ލZϒ�{�,���Z��cƒ�I��
�8$���v���-��$A[��O�N�6 %���d�T�x�T�R���ɇ���U�s�Cʥߴ�+7N���[�]�2�Rُ��C��v�9�I�
��םw�=�ê��W䃩��nǣH�\��-�3����}=\� .�n�QR��mB-��_��ɚ�Zd�2��Hf�0�������Z�k�$a�JG7
�?EΩ�v��;�0���}�O����Qaq�vr�!���KN����d�t�`�V�!A#�Q-��\�Yl��A�<����XL�6W�n&��bw�2a���Mz+�vP'o�X��"���Ҿ�FW
���/sCj�eo�5~�جCw���"ԴT����ܿ �b�K2�%5���/O��_�C!��΅L.�7�qhe���ď;��Äz��hB��V��	�5Z�%����nJ�44F�����N�wsS1`X(C�ãݙR���!#X�hH'rPQ�nOl'�Eƛ�����/la��_2�a���#��<��U�w�� �~wM5I�w2���Oѐp
QpP�T�<��q.ºGR��Q��+Z�Ԋ}�E�}����H��m�[oԩ<��ꡖM��me���^�̥�}dhԦ;a��\X���ZN���i�[3��	���#�Y���	���3�]ũM^��1�>������Eݕ\0�v��ײ�?�h�J�Ʋ)�B��	(9��Ѕ�*����Aq.��G4�'�6o�F����u���	��g+�;�P����������""���0TVw)��^=�@���y�K^����)��B��#(�<�w5�#����iGjە��a觫�<�΁q� �M��v�PE�������p4�"1$�.��؉�?7���Nf�`"V9�Y<�@�RY>.��m�P����< �kâ��~���bC�TY��}t���՛T�id$계<���>�L�����Ek7�A�������1#:��G�pog,j����"�Je���U�?Փiݹ�U�0
����cy�@��o!0��T���H�$�}��h�5^8�۷�kS-oX�,2|P?��+�t�S���G� �}�����#.^��ߢ���R�XkY�ih��2bU	���ʭ�6�fLD�,�v�
J��x����?��W�᫝�:/Hc�ۦ�a�wҶs}!��鱭��ҍ��s����M���+F�MK]�YH��b�̎I�^h_:
��hF���җϊ6+�r�r]=a����%�0���f/��ۺo����ڂ���������Rg��t�nCSI���u�kA8��I�:��;K'���wz�hlb��)�����6<>6���O�]��g��������{a������ISԤ]����L'j�h
E������V<U"N�����  Q�e��T�uyq���	��̸�e�oTe�$��t)�v���v�Y�ȹ�[&���R$zb}[Q?QG��N��RkEADgKӱ����ѻg{W�K�Q�u�Q���"{���!��3�~�.5��&���ƣi�n�k��bb��L�@��%�8�
��Mc��QչZ[�}��`�?.� HT��w�̛UeRq��z�=�ۺ5"W���'OT6CQ��KKW��%L�_[=���G�]�Z~`�`����X`�4�;>�z�������Ҿ����1dp�x�����L�6Ξ��אm�1j=C�8y�d��U)ĸ
��3ش��6�-s�֮�}�3{~}yɮ"��ߵ������!~�r�.6��~%�ku�n��(�^�c�����9A(�R��-`H?�UG��0$����oU��x����icX��#׭�I�ZN�����.,#@�	 7V��^Uq=��ޑ�&w��l��e���?�b�� ��<�&b���ʛ����*�"EGE wĳUVR�CQ������fѼXX�v���7�g�E��(n�e������'8[�F\G�*�3�KQ���%�Š�e|���!�z4+�)O�p��xaUM�X�]��D{$�S�ѕՓ�WOFL|'�3�t��������C��莘�.$;�:H�]�܎�m�����<![�MA�Τ�gj��7�N��1�s�b��ս��{
�����7@�F�1R��"�~+��;1+Fn���1*�f����p�v�[�u4# �3\�<R0�0y�a��d�O}y5��~����嵚����.�fa�������Y
[�/q�f��u�4��H~>(��9�j���*Da���,��IE=��Ǝ|���{"�4t.{� ��-�,t
���#�%��\�d����/)��q~����}�����
��`Ue��ug٠p�y�ܟ��n"#3[��֥7N&m8,)?݇��mg�ٜgy�&М���aH����������Qq�K&ſ�(x+w�'k�yT@!��fϼ�!E;�A"Q͊��jl	kl�P��3��4Y����k��Ew6]��BQ ��+q�OO������6*Jj_�˟�={lG/F�{��	���8.�Md��'M|���UP�U2���
�\#�	��%W��w��گ4��T��[t�����D�-~������R�ϒ��/!#S��_��tG��c(�qp��[�	+��}��y��d"��zϣ7{��/�c*�k��^ռ����ʑ��%pV�U��v��p�B�Dz����+���0y1���7O�os��%�K�=|�e�5�u��h�4-�J��a�d��cC~�d��g��}��a�k�鼷�6%+�<|�	>�0g������z��f�#��
y ���h�Z`q�0E�>
���s�\�5uQ�?���S����a3��d��J�"C�N��pk���������"�o=�j����Ӎ�w�~�B��κsIbI�` �d�) Hd�P�T�1b�0V4\�0T�[J��L�6:X��3z(Vc���E���H�JJ�}�M���nc?DCSpt��G4Dԓ����z�GL�A6��H�����1R���lp.d�����|)=����E�n��{T���R�x�{����A��ł��vN3���sOc�ԩ�W�靷q�l���ֿ��ʮ��q��u�j5��8�dv�]�@N���i��7�*�7V�H4I�-�r�DȊ���=5^��0�����<T��p&�#V��f��8`��X,k���d�6����5Z�T ^K:9>��s��~C1����ZU>�%e�w;%��c=C�$US���w��^��J'���;��tп���#��0��ccc�	숗#�_�c�-���ӧOe[㱉pQE�CҒ�J+��a�x"[���W�{�;v��G�ܑE�C@s�@q���1Q�n�!L��P��caaN��6�.���sb�a�Ӈ�rz����n ��jJ��hHh0��`��E�� ���LkR�~)F!��p��EL�ս��,;?����:>���yӽ�&�h� 18>�����N��Mv�'YH��j8LR�nWY�U{��i<���1d� D�j7뒗���,a�#.�3>���+`��9��L'7,9�D��z�2������,���c������d7E0r��:N��?4qΗ�5���D�D�8]�����[>����_��B%��5��	7�	�/���2'?�[�tR� d���� JqYfO��ng�tԳx�q-hX|=۪Zq)`�y��+V��kOz]�\LC�\���������xPֿ�5���Z-���;.��?V�r
#���;R�����qoŶ[��=����KLf�K?(�s����y����$_隇��C^@�'u�1���,�Mf�b��0����|	^N�� ����^�,ŐЖ?�3+��$�^�*U��渙�^Hk�]��q9;�F Bt�H+����4۰�YG	��X�p[O2�S����m�.�t�{m��b��?ã.��˾1���*�UJ����0ϧ���,�2�� ���3D� Rǯ!8��X�f.׋��iǴa7�������u�*z|�/�P�Tw˾}*��M|ƴ>IXي�l�"��z
��M�2�^	i�G���U�{�}���X(��e5m�����'��F��#s��3�e>���+��3��)u_V���W�R��*���@0<��
o8�v������oD gr�o#x�߄~�<!��NG���k|��w�xŐ�bkR�����5T{Aj�d�s�?�����Y����n��"��;��zO�-C��_�0�1�(������^�D�9�F�m���Os�"d_�g�����rE>���&�q!y���BW��觃��z-a�vC�;�@eK, "��4_kj��s¥�l�������6�<�gL�n�ߣs��Q+�A�\'���#��A�L��lb*����.CT��
eg|�3��|wrg`+us�Av��Z@9�{��1ji��Q�k��O�$l����V�ٯ�pʀ
��|
���	��{ec/ Jz����a(��D3ip�����a�Q���vS�clE�5���)����'ͬ�3�a�ܘ�X�JC��%1���)vf� ��&��~]����y�l�"){��K�Ck;}B��fހ,���\���y��l�DL�t��g�O���tl��@�F@��A�K���~$"�I�c��V7Qzv���ѥn�9K�Z4�¬	����XS�bu1ڱEJ�fK������������I�Å�%77����'�5�\Jg�z'�o���l�v��農�Y�\E�߈P���\�R[��*j��
�u��N���)�u\U�h��rb��dW=˩�>�W�z%$���^����y����/�AT��9�59�H��7�He��#B��=ܫ���CDF���M��{���|R������#mł�i?%�2A�e�r{��;N����繣֣ᢹyo�ӫ&���z��=�4s�:3�1�Y���㜚�q�j�H���)�I�b����HfÑ@�OK1uL^^����U���\�i�[���؏�x�p#��_���*A>�`����M�fԸ���� �YX���xU���1ـg�2???//�A�AA������qW��h�0���f����Oq��l�>늢U�Ht�k����Ʉ���V=�Ϻ�d-��Z�x�fc���阞�z�C55j��n�Ӏ�ĵM!M�K��$�Fe����ּ�[��Aw�.D��r��n��q��C��7���\��὘��T\��|�W���:M�G��V���w�&W�:�nD�ޯ�]W���f�m�j����^՚�:i��ω��=�X-��5?Sgcl(1��X^�N��.>��ͯk����������D\j��f�5x�3�#,OqQ��"���[L����X��*�!5�[v`�H�a��
��?��WpM,q�cMy��el�_��b���$Hx�$}�p>-�!}wOJ�aXRR�=dt���U�����8�ʨ����@ ����	��w'�[p����{pwww/��a��~ך^�=�|���Quέs�~d�}�Ѧ�����f��@Ƭ�%L�K�;tqU�Qw6������V8YT�wH����灩���!Cf�6E#�d>Ϳ[�w��a²Ju��;F�L�Re�=�>���BbHs���Q`m�Q� $=�V��TGV���0cr�)rV�#���9�K�w��h�,�xf��uZ�֥�}����#����˶������sZ�ظL������e���)�ە��Z'σ�2T��73�V��N��>
���ȵ�7$(ӵ�wZ��/&h��6���{�`
*� �����\]NB����X��K����T�)�Y�%�����1�<�i�xQ+�J�}l��(R����,���j���l�c.0��E�Q��<��f��F"�͜<�rz<�`.X�����S���Zt�|��[��Lϰ��u�6GO��O�C.r�0��"�P"u � �彠 ��إ���LrU�r�MN��V�J� �UC�a?�tg	�_��YӚ~[Y'���,��ϣ0�ξ������%S,��Șj�4>j�MM)�h�$�c���=�V�Dk��~E�E�������lF�^cZD�Ј�dw���ӱ+A��".yaW���#�MS!��-q�CW@�,R�ICL��z�˛��UP$&V1׋��4��,�]ӽ�M-�d��j&�q�#�D8C�c��,�����]�\N�����t��+X�5ůp�Ci����p�>h�.���6>~f���Z��@L�,\:�H�+C� ����9����� ��.���~��	3�"�kG�T���ַb]�ᶱa���+;����h��S�E4уؙL�}*Y:�O[��+��ɧ��Hp[ݗ�$���>{�2>;������ҫ׏��+�k�{����0�v��I_��l4$H
���'��5Κ�E���a`��U)UC͛霃�_��|6�J>���Z�[\�U���5�珘�l݇^�?"�I�yp�m��'��|��Zr�{��x~Y��)B+�������^/�R�����faP�`�>;f�+�U�9Qw���+_��3�wwT�ԟA�y�.�d�%�^?^��>��}�T.���.�Mx��E	����8g����m���;�K@���x�3�w��]l8C��~!����U}1�*�G~��n�~�k�Rr������t�w;�|���/$�7����$�f7T��Ma``��Z��n��!7.�$����Z1����]����q�Hߏ% $�$���iz�ނt&U�D@����2l���P'E11r/M��f�04NA@!-W�[6�._$⋮�E��b�_s�w�-����O �����(竀�&l�؋��ٜ�S��Hw=��ߩ���-�@�~z�9pS�`���q�''2dΊ�U� 1�}�1���)�u	�a/Fy�X�c!M!�mm�q�l��j$�aJKK�~-�{�7C� &3����:�%���
t)W���~E��]�@�P��a���	OS�<����%�淥��miF�c�����~P2*?S\a_7k��K՗�C�(8�&���#YB���;�K��_����5AVh�.�FU�?W �
SZ-�������mB�8 ��C� �L�������G�zzB�˸��P�h��P�_V��1���hl����&E��X�\t��:�-@,�(���T�r��I]Ҋ��S��t�����eƈ�h:�ǔ�+�8㜰R&Փ��][?'�����W�wC��xrq��������&}#ܡ���g`�y�U�����--8FJr�Un\ܿ㖪��:Q�x�Ʋlw{��%��b�%�5˛W���2h}r�l|Ӎ�MQ�=�]������I��yY�J�l������[������ߞ�"�����Y��;�,V�������jXb�x��Lw��?\H#�+ַMԁbH|�7+�y_v��!���F�Ӏy�+:&�Fk�:��}x|W�'���y6���ۭ���ɬt���(�Se����`-C��%�2�+����?���E����p����]���YCj�q �q��xA!Q���X���2��iE$;�9�v�z�HLCe�"-G?Os����GX{1U�IVQNt�y�8�F�{ӟs�<֔���m�1Cym��!o�>�ݜΛ0���<�^�|�����o�-,���q>:����kW�'J>o?"pl����2��sG�B!j��דV����%�f�&��q4`���Q��#.��0Ь|��(\f%��aW�s�?����\�;l�~S{�y��)���jl+z���<_r�*�D#V�$l����P�x��h��R.xp���i�;|�G����O����=��s������j�S���ЫJ/�Ԉ�@)9V3U�=�/ΈH+�1g7�m�7"���c쳛e�ж��E��1�X`��鶚K-?;�����i�&M��pX���"-gIqF]嚵���u�y�?Q\`��X�j6u�?�Q;A��F>��P�eb��|�E�|>���m��S^�vj=��u��0��h�H27�'���2����r� Q"����ve�\�h����-ؑ�7���
V�^-�&�K�巶��BR�l&����������r�	kb�#k����3���x���6b�k�Ξ�n?���A���Ϸ��t����#C��#1qpR��n�>�wa��o������ȏY�W�ጕ��[�]���can4�{����'-������*��҂��踲��t����s�;-2�:lXzB�V���bP�H����[u�a�׏�g�	��z�0�����a ���0Pe�������f=�l��4�^%�r$�p|��!�7�
q�����ǔ��&42z1�a�gN2Β�%ʹU���AO�D���S�0w�~$�f���s)���4۩Ef�����أۋ��d�9��^$�Pȕ��YD�;�]�W�kAz`���0��Қ^��CL m5h �V����F�l�(h-U#g�,bGV<ݐؕbeR7k#H��@ZBQ�b����1 m��Ll�6Qx�Ѕ?��g����7f�:9E{�$���ێ�}�y�&�B�"��M��zL�_�Q�bL(}�9�͌=��\3�O2��m��᜻	��Z���O������ S24�^�%���[l�J7"/cy�XN,�`�қ�n7��CҜk|8��?�!<�OGtP���8��Zi
:���yܐ�3��J����u���x�'�8�&;CT�P,�y���
/�wЖ�yG�YDW	�=���Q���G$��W���2�vT�DPqG����C�JX�$��#.җ=���
6�`�'9��}@�ܑK;���֓���>*�׊������ûb;����>�5 y�[�y�༭\C��O��&��;h@Ț�Ia�A��5Q��c  Db�J�״�0�_�<R�-��d���id}w8{�ՙᘻ�(ޢ��$�	�K�б��=��弅��y�?�Y��8�9����`������.Ŏb)�)
u��m�>ՈF��i�X7�c�c��˭�-�Vvd�S���4M��wȒg1�F�K�:�����셔��+O�f��}�����B:��j��M�+��S�{���{��o��ky�+'P#��[�����"����9�֍
,��f=��!�ROa���UG�����ci2c/��{H7��=�t;�*<)���OS��k�hp��5�W��"��1�Æ�BY�tc^y3��v�y�s���<���l��U��wΜ�p�>��\�+���3�)�k��AG����uwv����'�T�����O4���Ah��~��-xw��z�<!���q1�A��>�W���?����k�W)��v������b炰]��Tp!<!Y���:�}�Q�Pxl�~J�bR#b�-h�p^G͜t��К�y�P.�-�>��պ�o�����U�ˢ�ux0S����_�r:ÿNL ��g�bκ�#Qqsc��H�Y~�8��ㆧ�HO�����ŌB���,�&�3�DC�"�մ��� ȩ!J������t|{�0^�]����/bO\��Ps��tFj\�}�̭MoD3=��D��P�y�k����%���-��`m~��Y�cY�UFI��1G���tF�0	Zm�+�C�3�.;Y��v������)����lAp��֦_�ي�ǫ�Y��\�N[�l��_(pKp�X:�D!���[��fp�V�>B#��\s,��eBs�i��!�gDϨ7� �(���s4�ס����R/4O�O��*�MdK�S8�$G�h����RSI�"wr
en�1�?��뾪E�V�L1�ǈ}�x ��D��c`5�r�6|+'�040&֜QK�QrSd�nT�ᠵ$5ȹ��g_B�T��l�b�b�y��oe�t�C@Q�U�妪�!a��<`�
f���<3����ђ�T�h$0V���`��7y���\P�(!�c^���<�
k��VZQ�mm�5�M���ѮyC��a���;f������=y! �:�;4e	�'�ܿK�$�T��x�w��T(�������R#�C��D\�&4�
��#��_`Q�����7$0|�Ȃ`��y�Ntk���iO�d,
����a�_�*~��d��0�������u�}p��:�����z�E߭��-�D�5p5�sѧRԑ\�O ���/������f�"�=�ӡ�Fz}i�Q��wk
qj�����z��V��q��ᤡU�ɷ���of�7��o�i�.d�(��rĘ��1��1�ͤ��̞hjwTЮm�d<¯~k1�h�z��$k�nF&X}���;��l�(�S���ެ��U�\��p⽐��d���3��Z,�Hko`���2�W�$^3|�t�qx���EK�%^�;�����ژ3��<��U��Qa4ހ�^� %,l3_����E߰B�t[ WND3|�D�����:t����>��x=/4�<�=�٫�B2;78�������fcbP���bO1������//�L�CY��w�a�������>S��8H�����R8�|��77�gC"�48��7Ctܞ�v��ئ����,}��^��M����ш�����r���<+5?���M7�����@����l���7D$XT���Z6F �$��C-��)cK��/�!3�x*��:;���#��C�n�4�(��"������X%��ZY�E��p��3fŷd�ftG��Y>7�	�ق6 M*��vORkdI�%&+W�#����;մ�N�߭��e?��ߜ��yJ�%M#ѥ�q����Vc����Z��R�p��_����l}��^��H3jp�x�u5(LT=��^���i��ri]�!�2���5�RV�ŵ1�QM<N���� �s2��劋�!SV8`j�҂S-ISul9��Bt�\�����L�Z�u��/�J`���j��ш�e�a��)o~$��z�8,&�1�
	�ꎆ�Ľ�0nߡ9�ԤzIz�,�ӈKQIDЫZ
&��R|>����!��k���E E����2�(q�Q9�Q O_Jt'Qˤ9r��h\O�Aa����*T�lEn ]HUW��۳�M��F�uCQÄ�oO�z�8��W~�>,֥t������B�Nw�dR��9�l\Ng|w��M�9�������lG�/�?[�w�[�52�y���a�n�K��A��\�/��OJ���wX�WA�6֝��S�W~xX���l%Ր����]�s,����t��D�q:q=f��m����t\�Ng�dD2o�O=]�@�Go��4����KaE�T|�1S5To0���,�/I����J�G�Z�(�Į+i��7�R����+�1��J~T�9�~^'&j�2���!j-��/� GΖZ\��%�Hf���в|^b�y�{�n��j�'T�I���O�~,�P:g�+ǔ����}�Ak�������f����N4���1G���5o��1A���Jkٌ9m���+M�f4t�Tx������B��J[�}�����V�W���}`0���������S��K{O%���x�iJ���|'Ekڢ~�S���k��
��ݷ�(Ua�6��l�uY��$Hd��?�C�T����yq*�]����⮸�a��I���Y��OE�e���h@˾��i�ڼ��S��!h�_�C�ȑ'(귵?0V�����K���p��z䣘U�Q���R��`�����"�On�ˣ��x�v.~�h�Ąc�J����.^;��s�o��tC��|&S�7����8�A��X�Ԃ���6��^;ݪ�߱���`���}ZD�\?8UdjY��y�GZ��n٫L{��˕�q��D�u��Q"��\�(�&�1��Z��z��%�V�ѤAۈ��'V�J_М��~r�V�4�j����T��j��ˠr\�Yy>�Ά��%?�С�:��j��蝄�`*� '���S�Q_�*�H�qb�A��MR�/T�m�ՠ����R#���H;��"��Q���(:��8L{����}�d�T�f������9JV�m'�U�
�>�~���V�ϥ�lw�K����F�;(z�ܣQA��H�����l������^�� ��Q]Z
��~�fT���ޔz���ڤ=�`Vk�l���sG2����K�m�/�a���v����OI�p8hy�h�5X	���yޛrc5��(�qɻ��2c�e�
SV����<�+|z��N����W�C\c�����P��۹�'�����7��Wک��u,�����l�N꿫��읠!C.��=[�N5h�_t:%�;uzb:'[��JuI�3�VE�黿�Z �}-aK��@+ܞ���Oo�sɻ|���}Z;�5�T����À|�ә����|�1w�V�[	�x��c��>�EL�����j�۷_�N~���ȼ֚�q�{QWY�Z����[Ezϱ�'�0�_�C,aFeA���K;�����XZ�6�KȒR��kU��鱾�~n�6�n�,YI�qǸ� 3��̲��7*DM^?�e~��U�_�ڜ��4M��0hcV!�>��"�~�!o�u}�הĸE��G�s;���vf&&�ڹ�v���%�����%�gl,�4fK��c���(%*����c���
�B骧o�0�I��QP �s�
��6[��x�qmk�Ӗ�c�r�Ճ�Wf�]?��Ӑ(�����ȃ�8I�<:�x�|ɼ��9,!�L&���c�:u�3�ha_4}�2���G��PWW���I�� |C�Ϩ�ň��_^[�9n3�����g��ᵉ�ߧ+���w�'Di�3�����f�H)�V�0��� kM�y3��5W+�I�x��?�W�D:�v�������P�]��T#�k�[mg@>	g�$���甤d� �7'h���|r�2�*��o4�N��NU�;�_.O�4aaz|(��i⤐1����w�G��%S��G�9�T���G��w��m�����u��`���^���}��V��� SM>k6� B�Ɓ��xcJQR��&� .��+;�'�����00��׊W1e:O���"�C����<D�\���lM~���%;x�DKot�;�W�w[��*iL)����ƒ�f��.��hiX��4�{��΄��L̯xJ�Z2�^sIC�Ͱ�V�P����p�vwo�a��*���ǮZb.2 ����] ��϶�9d��x���`��P*���W��a`���n��9z�9Q%�H�Yۑ�^$���w��|\`ш'O����N��[ܯ��q�7�%�0yF\���_W߯M��F:��Sb�N�]�v��LC�iѡ|}e�,���_����f*��r��m�;7c�Z$}o������Mg����вk#f,ɔі�o���� �uM��YYm��M��n	.�~c�f���H�jb��WtT�@��K�H�^���*anY�ESJ�h�L��z�%�I����`ZN�w�@j,���֘^��-T�����V�WG���N��_�/�|hXT�z�-�ZK���S � xYz�F��ܯ�9�h�tj�������vU�(�5��{�Y�������w��X��1�㢓$�˵	A/~Z��?�&�_�zx�3��t Y�`�D؆LѮk�U��� ^�(b���Ck�����T��>�?{`m)�g4���3��4Pc�"����H}�bWM�3Zs���gx�5p�bCh���J��[��%���㑊?��Ɨ�ۣ�Dg����2��Fˬ�S����+�ne��:>��3rYhcrT"d����g��7���[���n���5D!`U�� OZ~=qŷB8]ք��S���m�&T�U�ؗ�| �Dy��l��[��ҫ���{ �ui�yA�KZ�����K*��Ŀ7�#��`q{w��x�r{�h����l~�PQ�l�;�J�\���*!��8�N�i�7�b�{��0���P��H˃��
�����O��k���LI2�ބ��&O�R=�?��BW���I���;X'�7�<��3�U�����Pɬ��kr{�+R�Q�"7Â�B�J�[��Lp���O�6 �}�Xs\Fp�uʧtS�`��dT�9<�h "�}T�ҳ�o4x���$�\��]��Ҕ�M'���d�ݏ96�'I�r'��{�T��)
7}�A�]�_� �	�t:����5k��P˕  nZ�U2����3%F��˴\ɻX�R�`L��.�~o2O�Z�T�}�D�b�Fh�ŝ����rw�m�Z��p�'���b��$������,E�.�?aC	���g䟧T�&]�Q�V�W�/��2&i2KZp)أtB���N���5p�2�rT�'u���;�K����6�7D�Uf h�K��wb� !��ˏ���� ͮ���r��l�$/�?��
;��oaXieEר��jr:l�)c����J����r�ћ͞h�L�Z��Z_?�.�;` �)�:�:���Ԧ��荶#��_=�Rmq$����g
;%�z��	t=ymX�<�rr� �u=s�[�U76��H5���.�U�����Uۄ�������M�r,����Tgn��`�BK��&x�pc86�1�.kl��:�it��2Q�#(�[`^Y�rd���uI@6���w��g<EDQ��7�1��%�B \�=�5���w-��V��,���|���S�z�{�NyE��u;�H\�W�����f{�{0�+
�.��E��P�'ф���F��)��[#�y��h�V9����p���c���%t��vtrz����0��0�;��� ���8�L4��@��j
4�hZ\KXn����]}>3�xX{����5g ? �e��H�!��*i���J^�������k��3Ol��3o���3���	/{x��VY����G��5LPe)�h.�^ �lz�sx^Y:5D�oi�T A�	±�	�����rt�$8C[��D��r 2��#M���^��(���r>_�
BQ�� �nll@���mm#*++���V���&�������<!��2��d�i����&��z`�Hl�c�y�AT|~b3qC�.d�WT�`����8��~ �9abI1i��i�6t��ݪ��;[��S!rXq���w5}� o�!���#ɍ+��@OO�6�7@"~� ]����D$m�;�R��N�qwEG����6RQA�M5�l	�Bc��hf��L�����h�q���$����b�Jt�R�O��l�G��_��3�+fR�����(E��XJ�1�Y#��7D����"��g�K���tCa}�����OÕd��A��/��2)�	z=YX*�&��t�F1]�a�6�dٍ�@|V���nwÉ.�Ԡ'N�`?�~�.K��[J��P�KM�k�_!����K��@vѵ�_�@b����_j1����xp�
��p��gSZ{�=�'~�$��Ƴت2�B-���xZ�C�
�0�ȝ���ہ�%ηe6Z�-B�Y�O�>�R�gg݅���܊��+�E!Á��e�2���W���1\��xWgdW�K/��H�_Q�^LGs�� �G<%��/�j�ب$d���]i�/�FS�My��%�3���^%��Q v�!X}g�<�v�������f؜�D�7^)	�K��1M���ZC��jC��iC-�h˽�[�y�� r�ߞ�/(�+ף����öa� �2�j&zL�2$��~�7w��J��V���
_6��Y��,<��`��)���G���f_�,��J������h�<����B0>Q:�S�$��
�Alz[|�>.p1E����� ����q��	Ks��TD3�b�����Gt=��`����b�Z�y�(���qY�R�B-0�h��9��0Ci+?a�^_�Q[�[���p?F��qj �s�I�g��i�٫ۋ���C���;`G���8�j�:�/��I�b��q���ҋ��@��5ňZ=M�T�4�-`���F��<I���D�%�y!Pn��n�7���㩩�ubG)�t���зYQY��(l�E��M�C���(X~2��bY��]����s�|�A&6��V�~p"�!z@�!^����튙��j�;5��Q��_Ƅ��6�����X���"�����S�pAL�9>q�����;��`��q^�QV�<�� �6���3Lb@��<w�c��aɡ�(�
F�� ��~��?Q���`}k����m<�0?�I(FQ҇W{�ꥉ�Y,:̽ CY�7��S><'��waI`��u>�0�©ݔp`��m�Vr��7i�]����J��J {���:�M|��g��pw |�VOA`��^YU�?���Д;h��AJ�s>.Θ�� �{��-���x��t�g�J,>Yh)��v4�?�Β(��-<W�%���T�@ ��c��+N2�qPx��*�N����B��C�T�+�D>@'8,3QW1Є'p/-��#}H/$��;*gG?vFm�|��/�����񄇇G��I�q�9(F[{{��Ƈ�fz�?�"� {���Μ�����$���xé�������h��ϛ2��J<qh�[���ɬ+n���׊@�����7�M�W�S��e��A�Vf�%A�O����v�[��������$��TʉzN�"�agyx߿S����ZOλEr�w��+3�?e�H�5ҟ�9�8�O.*ܦ�v1.���
|wp]�֯����4�������Fm1
P���!Eƙu�s����Ҥ1CYT�;C֔ ZK՟ˁ3��.�Qۊ~&5�B���_��a!���\����a/��H8&5���3a-�,�̓�U[w� !-�Ggw��L��cv��'�ѥ���������-,u�m���c3�t�&ْ�l��r4Vt���o�B56_R���<�"{���4���D\i�K�~��!,È
���s}��2H��t� ��+R���_6����N�q��W�!$P�@��H�
pT��V�Ds�TC��'J	���.R]7,�p$��h���bâ��J�W�T�Mgg�<Q}.y��"�]m��[���>ͣ�nR��,v��]���\�-�)�Q{)�Ry\�L�v�#��W��T��@P��
��ih;���.I��؋�(K�U�5M�S0���ӓ�ѧ����'��n������Tѕ�c�R���o-�|h})l��mm|�G?���444x[E1C�����E���� I�X]�c��F`T�����5�3[Om�}��*�Mj�홠o?i���K�Κ�̏J)A��#o���r�ߟ��;�S�H^Cm��чM���6�7�.��d6���%�ū��R�G_M?��L��,��U�,�ކ4���v�.�a��MAl|C���VK%W&��8NB�/:��w]n��������z�3�4�����.�b�@Ոj3g-YUhK�TVt
�����W�no��L�d~1q� F��~6>{O��V��Nw���Q]g��"��"j�H�J ja����j����K�-OàF���=覆����I8T�H.��Gq�N[H䧓	�*�aG��Lzz����i�"	�{T�O������tP\"��y��W��Q*����g�J�f�d6G���P
�U�ʨĲu�F��N	�Ƞ��LB�x���Sb*^�e�I�)'�G.���6�����Z/�*���OW�,�������+�Lma�)��q{���[vt�5\U�bY��b�����Z���.J3H^c�c����t�zr��If=!I��������g�%i;�������/��hna��K:�듩���t�����~�_�gNΔ�F��w����i����B�߼׆�t�w}�(�3����H]�@���y�P-'`�<�2enxAU����Ϩ$���Q'	v�ihǬb��ӷ�����6;~T����>�����Y���ͯiP�CL� U77����_2(�&��c���>�pFz������/IĸY���d��p�/�(�]1'bZ��lZ�M��YlEj��3�^	�G�}�~~�w����W�?ZB�}�V�G�BoȒ�sAWL,�+q���f�����ӄ*���2|h>� ���Ѱ'���gh'.��"Z�z.Y�:��q�A2P �=$�u@bi0;DFv�"�~���'���|ׄ��C(��]��N��?w���&��0��:xpO�{7�Úb��4p��`�ɤ7=�.��l�\g?G��pBg[<_��b!��Y��옽1,��C��g��tv��}��~�����qq�p;����!*���z�vC�(��W#�)_�IS���9�ly���Mi��W�[�����x*~pu�0���è���"��DDH�P�X��N��D$|�'������(n�������?�����7����fI$,�{4{]TzD���e��{�4��)�����M�%k�?N&t��6-M˧pͫf��ܻ�I��.��5�9>EB�}���N���9,zN`�� ����<��������.�\�KCڗ���m�����H@�z���|��ĒfǱU��n.`�0�S�Z��;����y�>�F-�'�pɻk�E�;��m��n�A7Z������P3K��0�ػԑ9�w0����������X�҈�T�l���l�z���>�)/�w�d 6�D�ql������&�cG�'a�B]�mJ�����8.)Dm�P�:�|ɔ����r���G}�\�@*�j�1���,�թ��$�1ნ/�?�79eJ�ƯE�������v�`�$��/+
��S�֯���9�4�5�4���aT��,��}��=��	!!�Q
	�4Fm�m�H��3 �C֖$xs��)oj�显���:k2���+!j��T*B�
6��-�X�k��<
O'f�Y��K�Fޝ�4�t�e|qo�gG��b	6^��XU�Y^�׽�lo��F��EQ��P2�����l#;d���(�6�b�5��e��eo(Gq5�Uv���w}Ol8�g
C��ep^��霑06�@%Gu��߽b �F��h���3�x�4z����a��f�$�����U�sd�Ι"�pG1Ĵ���K�����jd�UU=[=p
����6c%����;�(��o��m��[v�ף���[v�W�.�: a�k�E��?m8@��W-�(��F6C��ݧ����m�R)ά��T�N(�+	���
��������[e>��Clߗ��������A<[h��c�$���`ɵÖ�F ������g�%��U�¿؝:�:��Px�߁���p:��}��L�����#����� 0X�����ܥ�eߣ�`�Y��:G5�p@��3�1y/���YB�:��׸f�S˾ȕ5-L,��}>���Q�,�B�;ѿ����6V�#�a ��"~��w��p��Diu����b~[3��m����G�`^7����Ac���,���s��\���}L���s���|mfR]v��4�>�m�����7?y�<8g��Fy�K)v
6Xc�B�d�R���'�Pi�q{p�'������|Iisw˄蘝�M7�ŷQ~0����Y;�}n��Xqw��
�Q�0��r�8�o9�5�á���F�<��>3D���
�-Ka-<0�!G��oC�����0�Ƥ��(ٹ;�Xdo��VWE��ZQȔ����[��&5���md���J~	��귒�����	G�@ˇd�f�S�I����1(�V�tȁ%�.��T�"(Q�;��#��,��s��n�lum�f��E�	��a2X��1I_4Ӛ�9xъ�>xvR��"�-����.��QW�{�U����V1��F�]�������H@fTƬ�U3�aV��#z=���b��tS��ۈ\�3e���+7D��9{ߺ�Q��|���0�^�u��af����v~`�8��Ias�W����aYʾ�v��H�Q��m��&h�ɖ���^У3K�p�fr�����v����{���.��v�0�Vd���,�(�q�Ϩ�ģ��P���_�Sև2Y�7���#�S�=M\Gyͨ�j�L�)ڜ�q�-�c�5~��x�A��&�s&�?
�cGSvFu�t�|mJ�mAC�}ڹf~�͊`ry0�hm6�>]��*V0z�A���򕗵��'��`��V	�6p`��=J>�n�3�G`���w��K�2O 5�]Y���hr�	�h�豱��`���\G���5�,⫼�DC�IP�]K����T�}��U{�pU8Ma�Jv6 OdH��
"c���[��� ZO��|LZ�������%y�+�l�˃PK��	f�ןl`�B�S�����{�Ⲍ� ���H!�m�y��,���1w��3t}/����m�(�@�03������g�R���@˨�&%�4�zi�C~-ib�ɡ�û�A�Ҟs��O�V��q��?�Qb�����5E#��1��)L��%@�%7M6�h]o��&�Ϟ�q/�ģ1���_+W�h@�cW���	:��!���}9���F
�̶Y~*�OoTT���8{���"=�bI�H���*B���AO��T._�g�Z~�^�)�̣�0j���b�.�=P������I��� ��&��\�%����Ptώ�Aw����ĿK� �O�d+)c��uyT����7�4�<\_E�[����M��������J���b:��!P��h�g�%�[6�e6@9�����*R�7��=�yR ��忊�lx���/{ ����i$G7!6����SD+��o�:Q�����d��
�h�fW�W���5Y�<�k����W�S��m	�V�$�r}�-c�j -F,t��:�kp��U��6#vpf׎k��M
4�^NGГ&,���/�t�-�.�)a�=oy/N(^CP��X�Jtޥ�w��=�'��`�-��:����8.+٨iUt0m�8���v9K.����k�e�2V��{�/�Y��I[�%/���t��Q8"2jh�FI_V�4�(z���#�~�OR����=]���r|$J	qL�p��usu}���~c3D��o��]�2L��������d�RRz^W�j\��i=�+�t�8�+�L�m��N����FY!I�s�A�,�rp��f].�]���9OWy����� ���s���o<��/>ίe|<��>�zy��(�;�%�X���-���A�H�$63XT���$�_�19&�@ٞn*�!��dep.�vݽxpMg�o^[���^d��i���=�g_��WVG5�pDX������?Y��Ud�����-���Ű����lf:*�XA�"�7�!kZVQoIm�B�'R��)�^C�\��'��7��"#��A�*�O!�ߎ�i�o=5�Զ{�#�j9Y���.��K��O��m��#~HX�mWTJ!z�IFľM�V�My�@��v)^�_�� \��̃���kqId+
�e3f
�E�m4�ރ��������4k�L�懃Q={j�.��z ��+��$��dw�8�^ڤ���e�I�f�q&K�~Wh.K,��G깾_ka[	�����g+���0��l�^�τ�B�M��u���tL����8��d���[Ӕ,�?vXM�D�1I�k�:�&��
S�(�t����m<�IW����h�V���J��x�D�,�L%N�Zr?_�`2ب,#k�cqw�݄����k�z�d����z�LQo8�qe��Pr��3���j"]v����"D�"�Af���$���'�$<s�3����/e��kO(1�G)��Q8�UK_�I�5�u}K���)���=���.a��K�c�B�6(�/��i("���r�������	����'=,޿,|�vC���1��LJ�4s02�7Y�!Dei^���3��l�s�A���i*�t�nJ�^����l�+H��bp�����H_�뻆�ؒﱸly,o�VEn�k"|p	</�e����?)O*�z�
�s�kLJ3��׷w/�<`���b��9�C���7�g�_�"��H&�}��ݜk�����:ִ�_�~3�jf3Bye��	�#���{�]Y|E?Kd^�Z>�Ȼy #���[X�ۡ{Qסr���m\�TIS����f��N�ߏ�B�t~����09�^K<�8E���I37�s!�x3?� 㱿5���$D(�UĒD)#��@Y���/�����GiNc�H�ȯ�TcRB�r�#yIoO<�h4) @'�g�~����W��r[v��G����?�pܔd���똆�Yt�6��/;�<U�����!@�/�[�����u��a'�����;��ު0��b1Ӿ!�d1G�xe0I�������d���1��H���x�[��Ҳ��+l��CJ����7?�;��[/1�R�k�^�ڈ���������޿DDD$����.��A��Q�nTr膁�`�������x��w��~����\s��s�u݋}���zO�ך�}I˝�ׄq{�&@\kT_?U��Ai\ی&T)m
������Ү��p�7O1���+�g���
��G��0^��r��@��eY��E�����H�;�(��J��Wq�Un(�l ,���%;U��ַd��Ш�$�5�Ml��#���I@�i�'�]�@�0��%��ft�8������^z<�W��.��z!�-T2���#�
��P���ڒ.�%o}u�s�\�Y3[�F����1����#�Z�yM�އ��υ���CLVg��FS?k����b�F��޹)���J�[�gfFt��r����8��L_&�~su`<z��3��{H�F�-;�J0~"��{��q�d�V��'� ���=��o|U�"��	���ea�ɭO9�?���J1�fjXhC��'�/���Y�;�g��
q�.\�m����w /���Ԣg�`}��ad�&ߝt�2&��ۆN�^~��ղ�k��MO��\���@�r���8*��l��V�y�����c�c�B�F6/l��~G�à�h����X�qta����4Ve���K�C��Y�;�y���2�5�@[�Z7��=U_���˶��%	���������A�J�!C��Cg-���y��G�P��E!Jm���3��a�3I��|BI��Z�&$�Y�o�x
�T���Õ��������Z��G�)�
�j�r�4o��5�t�_���~Z+#���v�I�y��S�r{Y��7"J�bU����&�Yc��)F�j��񇧞=9��+�W�=�p�iЬ�fY>�"s��>3QL~�7�� ����g�J�>@��W��m�8�TT�`��j��Ҳ�lOƻ�v�������/�qv�=Q��U��Sc���ό�I�}�k�w�t_�0���� 2�Q��W�h�k�=��n�0B�)Aa��B$�� Z�l������D�j�3#xi�q��V+��LU�Ic:�a��}���v��/7��Z�s�~�W��)�����ٷ(a��O���r���72uO˵��y��\ބ��Cf��������H�)K�᳑��h����F�aZł������k�iZPI(�,��=�՟��* l��wD^��݉	��Đ��o��_���ӯ2���^ӿS���{W��w�\�`�����dG��˸��BVF��O�AJ�9ŇݍX��= cz�1��&O�s0"������)-I'�悇S��~y�XP���39���ptk\4&�Y�@�'\�}�u�c7�巳b���"u��`�,z�'���Z�(�]�;̀�hܞ�8"F�����]>�#M�ȌhtН�+��i��w4���������]E��r�t��a��^nel�m{��o��VE5>�f]����?��Oh^��f�}�=��d�e�������ٴ��{�"�eS�¸#=�l�ϯqK$�j���� ����'�~B�5w�^��@�"��>~���t��DkM�Z*��e�9��B�SB�Nl(����8xb��<�{+����y��w=��:���8�I`1��բ`o�����$ȏr�$Ii�1�k���7-��(X}�"QH�Y�f�U�m��oFH���ӧ���m	2x��y�UQ)�<Yw"r����9*��6Koj�8.�Y;��A%���#�@�a���"��,H���ËըJ ��I9|�lqq� R7�O�+�ԍ{JO���c�K�2�]�uqЮ���3�:����7i4oW6=��%�9��+yk����I����������";M<�qV���dC�J֯c}���F�~�J�D�WF3\c�\O�rÙM� �b�
���p%?��u>^݊ݘ+���;����r/�2�Gw6�"n�Ef��=&���)���M~cάۮ���e����l˺��C�vm�/��\F��OVk�}�
�����'��j�M�}k $u�8�����9(���T��
��`�'q�*����B�'�Y�jNe��]Y�ʶ�	O�'O��'I� "ZUV��"�dLb�*��B�х��������q�ߊ�sD��jrS���	L1(=i�Ia��5�/�J�ړyt̰�Oթ!��~=��������s)���[�w'��gU��M�ߕh[���ieՑ�Z��2�r�y���b[g���� ���>=���k����Σ!���ϱ(~񟴽��,�c/��b�ʯf7Eh�.I��6�������[kJ
I�C\�o�����+�}����?�_`M��GO�|�K����/���"ߢ$�E�Z����� ��Ug`L7�~�
���~��o�.��9�J�\�	��z�,bp`E�^ܚ�̵b��P���P��T�cPe#۱����\��^n��g�W�Z��X���?8B��P�{��$6<�SoH�Q"���Ƶ�7E'�g�jl<I+l>?�p��U�e�0l��.���e_���gH=�J�y���w'�����$���T������d?�ůj1G�)��8�ds���f��gtJD��Hk\ɽ&�»ֺ�� ����h.J�B߬;�;����\#�U T^Ԥ0���>#dN��2/:\w�����p��׃u=�fk't-��I����/L2m��]t��:�V�(�*��p��K����cb�'�J/���B-�O(9����1u3RАJr�I�2��cIKx�KZ-�~��B�j�tt��?Y��v$q��	��̎1�t��M�� �F��ە�eR�aNho�E�ֶ���᫗P�1j��'��f���ȅ�?�����4+ݘ�~O
�
��~3/X�N���,juc�uj|e8�5�?k"]>�ͧ��x�N��3��)�q�]�]�37p��(9_�Z�om׻F�b��v����(�Y�Y��錳~y�Q>����@E�]v����6I7w���{�L�RQ1�=�9�.MAn�-�X�����~��<��`�)D���j��J�RU��p����A���G ���p��{�A�X���C%��P�a����.���\@�ҸأIJ��j8Di+Ms���]���*#�Z���S���fmptz"hp��m����y�QN���m$E�����՞�7g2l��}�#����Ak2�����z�����ߟ*�-Q��@~c�X���z�@��i7�֛f�����yڤ{��d�?W�$1v<��sp��X���=ۏ�y��;�g)Ϋ�m��(+/��L����E��](dd�a���?�U��D>�Uc��n`}�`�2���߬7��cu8�g��i��悷�JX/�U�P��(�������s���߭��N��YX�����-_�h:��S�j<Y��o��[�m7=cL�"��	ȍ /F����#}�a�򵱺��fI̎�6]0a?l��ˍ߯��A��������3.�~�lL�/U�^�k�kP.�����cx���/0fh'��	�=yt�\YM���Ia�$v{ ��e�i�|���:�<�I�!�`�E��dV��Y��nk��N��J�f��H�`Wמ���ĠZ����mZRg��QLE��hlfqi���QDz��V#������Aox���T嗎��}��t�%Ģ��r�n�vp�G4L%�>����DQG�oW���F�����m��i�.��E��E2r
���@�Ֆ4m-Rx���<�m�
�ݫ��6E��^�/_��~�#N9��dް��N�rjn�͈2�2�b�ڸq&�w���.��оoج�4�Mb�T�3}�"�ɂ���HrL�W���n��������̧�.�|^�x6�wO[2�J�^�|�sx��r�.I<.����	�N�P�AGŌ�+��wI��J`��VjF&c�E��s���{�^�~a�_�I?8> c��8m�\
&~Ⱥ�.aT�m�sWG����Fm���DH��;Uv� �\�7���tr��R�,f��mr�,�^ =��l�w�^���nD:DCGI�AƧ?�� �B��S*ݥ��U'�,�@*�^$��LfM�Մ�ǜq"�n�� Sߎ�_)t��>S`�y�8W�2�H�����A���7M4�˱8_�qB��ƮT2a�(�h�*�M��,����ȄEY�3B滃��TAf�d2ws3)���I��d�TSgV��Ys����)]U��D�@�7>����D��VùC�m'���1��(�ƥW3�a�i�G����r3�D^�G�Hb����E�v&ߨ�K�$Q~۲-'H����(�z��U�����=b����ѷ|�+��/���}#q!���#װ|#�P�r*�y̠�>Zd����v�g9��ػj��-H1c;�;l��v����ތ�C�Z�:�V�w���l(��=�f?+R���O�y�ٞ���S3����2�W����|�b�Y���˽I,�|Q��V���wS�v*�L�ඪdr�
5	�{����t�|h#�:���iʅ�����ݙ��4:��|I:n���6��&�W}�r�@�l�D�b����%(�$6�fs��|��k��b��4�D����~Sg�xm,�q1"U�W>��Qz'�,��u�!U�B�|���{e]N��p�SCwC\+������f���Ʊc���Q��;X9�ճL��aGRi�IޞLs&���P�emNd/��([�^���r�'�n�&aQ�%�W9Q����y�j��Ę'��(&�>�3Kg	<����* �����ИүW����GlƉ��p	��de(Z� ehr�������z�����QbXx�������+3#�[�q�]���u�8��L�$f�B�"��kE��(D/��>�zM�PUI~:�\C��R#�A�����V�C'6�+�x�+���ÒI����Y[���8��;�k[3:��J�����N�?������W��n�'����#20Ay�{��I�/�s�3���K����e7��yF�|�*;e�7���
h�L}��D�k��^7m�V\�� �)0.$k�mB9K�xV�{����1��%��U�N�A��
pϷ��SI:qqե�%i�S:�_�!��;Kt#�S�M\�<̣r|bZ"�(��W�շw]�7ʰK%���7S\B�jX�z��b�"	�;����}+�UV~7���o���g�]���p��{W�^[ۤWz�J,���r8�4̙��)\T�zA��H��>�r���m���������UG���w��\�ס2`��)4X�ϴ�tY�(����d9c��<�8٢,�Gq/ik92���zI�,u����ډ� }���L�G��=��Lei��*��xW�N��+��ݢ/��A=aN���R��o�?�G���Y�����'��'b̺��S����,�j�O��s�uX�wG��?�%���F�s����e)�e����`hD�����L^�a��D��?-����x(����!�ب�w#ef��P6#�Y� ���d��:u�Ƥx��5YL�*p>�G��ջ�ȧ�q��6u�SS��m�gnDM;�͘O�!@��*qP����F� ����ĝ��+�2c�B1�*vo��v�L+l�Z�e*I�RgF���!DhY���O�4L��I���2R�X�fZφgx�(��Va;K����o����}�D��Ν%�J~�/ ��Ы�����J��	�y5���:���K�/((@<���M�, j�?��6;�O��_s��9�M���fN���1#%~��Ϙb�A�,�:�^�a������K��{| }�@ sra���5�̺&�����}q��m�+}����r��~���W{}�*�ӿ�ҪGG��J�E$�L�R�'��"]��Nee�[|}�Z�gOE�J�3�$|����CZ�L�"�ܤ��d Mn360����
�@���4n��rQ��ɣ`}�)�ׇ�G�震}Ua�����.Sa�l��V��6{��ǻ<���Tjg���Z�_::z������9�L�{���Cw�m�����7A��#�`$|�
� �����w���,��o���@z�7]|%m�n�[��ⅿ�L�un��=�
K�q����s�!�������8��?7�Q���)í?B��|�_a�t>�����\���9�)���0��ۙS7Ƣ��A���i�59����iW�;|�>bs~��7u�L��Sr�$W9�����o[�C��a1�E�_S�z�'��U���`�%�gqϗ �������Uڛօli��|V��[2n��E\�Ьf�8d�؃���dQ�JG!b�c��0H�y��=��z%B�|��Nj'D�����V�ܖq^�NqypDl������(Ty����y��$���z�������$���C#�G��*�H�K=�/Ka���L�r)�p&��e|�<��o{����o^>���٦��Dl� 9��K��V���v٤������l�r/��0��5�D��w�(�L�O0�4�C�8��*��֎1�����jS0:*�x�>�na N��+UK6�}��1i~����RhgqJ���*1z���}����Hv��J�)�أФ
�1��"ʈ6h���ͦ�)���u�?�_�YdXJ����|K-�]|-,��o�'DZctSg�X=��g�x�J,۳&�	�WH�P<��Jp߮�/�	)%��8Ќ��~Ȏ�(��ٿ{�� �I��z{�b��N���J��@$ҡ8�SyxV��CjK��U"�nF�4������
S����eA�R����L��y:�m�ٙ��E`�.�b.v$JxF>w��eÖ��y��R~�wN�����Q��Ma���}�R/G���Ƽ� 9�ك��������F�80���r���K�+�B�>��V��A��m���eL��3B1�d�Qf?��!_��Կf���f��9�����9�N I�����\& S�8ɻ%�ku��1Y�"�d�`��7*D<�Nsߢ�;"���S`�f$J��&��)�v��*^*Zz�E,��Qڋ�d���5��
oy��l��V����Ӿ��@���U9\�Pe����-9��縮ue�XalK��]�w�O�zd�O<�U?�����h\GMj������8Ѧ@��SD���&\z�����F���.$�I5L�Ex���u���owb,�kn�q�U�@�(W�8}o�*��_�Mz������'R/ 6D�q�p�q�n�2�XiO:�g�U��f�e�r��/�zG(ǿ�Kʴ�.Dtu���tT<�l���8ve5�q	�@�#N�:�nq�爗�ߜk�O��0X_g�lݩ?�[:i��wѱ5�,+���P�����3Q��0���Lg� i�*d�A��\L��5x�� D���Kc�2to�c�o��`�� ��iD~��N��:�Ϋ����bT�O�d���;z�Y�v����Vj�x�W���&m�����Yͱ�G���� ݍ	�0��!�Ѭp%u�����`8x��夨��f�lUX>�sL�<%֎=�fQW2)�H`��P���z��ܲ߁�(U�)����?�z�`�F�`)��ul4@�ّ��B;�sx#���a��)��y��*�ts�I��2�t�(��,o"�Z�����,�t��3
����+;��AS��Y�s�9A���1NY��~4�m�eK]���Hw����G��n��d9�����~�_M�^�U*�]&a���Y���%�u�0�Ȉ���F7ݩ�e�qP���xߥ���Z�>����O������JT�V��,6������d����@�t�F�{ڲK��Qi/��Qǡ��<]�z�ق��.e�9��hJ���w_A5����(:~1}��{�m��Lw�o¾���E���[4xgerb�ǑѼ_>�ي2��5Q�/�2}Xƭ��1Ypز�]*��E�G���D�Mn�7R��)T�_�ê��=(�����˄��>�Lm2o�]�q�)BX����p��n~���N�n�n�O���1�qP�W�7S 
a�7��?�#��B]<���sw�q���G{�[����3y�#8����Vt<�R?�XC�=yl�m����֘���L����|������]4;���+���<�C��\e�p�NԹ�J'�o��>�k����ş,�{dt"1���ٽf@g������0��"��6kA<y�U/dg9<!�ٙ#`��a�ې��������2V a�9dG<��,e�� ̩�Q�|eԆ<�����)�"��h�����K��9��ȾQm}�j�b�Q�����'�ǯ���;���d�>�3�`����].ي|��K��oݘÕr�Sܿ�S\X �O��,�e���zRo��4;$�ר�(,����NL|/d�y!z�9X�H�ш�j��ss5���i�(M&ٟH�������B�z�%�wM�zl�}BqZ����J�8�[R�u��V{\��V�|��+��9A���I1]������Y�У�1����� ��K���ph�����$���4�p�m9V-���vخ���٢`�!�3u�����$�|���B�2SI�Ӵׄ�"���\�����5�ȉ*��.8R�֌��ӗ?��"�L�b���96w�C3'�̡q=Vc9T�ڤ���_e��s���剷B|X�򽺯d��By/���E �8k7{ z�qt캑�1�w�y��f+�Q;����ࠑG��!�������`�L�Ȗ�,2��+�h`���Q,�� �J��!{��@���C����C��D.��I=1���սCcl�gq*s���j�H�.[�`������)Zu�"g��k���]SJ���*t����5�ֽh,�;*D��}��{Nhs4u��;����q�'�p0����꩕�c���c�abi4��CB|>`m�����V@տAx���h�fhA(�B����k�g�@uH��d�4��ϛQ\u&X�:�\��AF�u;�)_gnXi��:v��$�(!?:8�����iH�G���^���u�i���[Bp��w&��#��!齁��"�o�%Upg��R�����mT`J����aP�Q1�C_d�ߖ���F�)ht�V�y�I:����^Ķ�xT��m������/ƺ�gv��c�E������]�!N+�li��c/��2z��vq��I;�R�Oa{L����5d��ơ8:��U�l�a�5J��E;�����.�a�X/[�*��h���CX�%&��
Q�Y��<e�tm�P��d��m�z�{m���j	�Y7��Q���Es��m��I�Y�z6�f���M�V��z��<4�^�`t��y45s��$-�W揑Ÿ�����9��{�M[���a�/��<^/LY
��[eА��sR5S1:˛�O�n���4�V��
N��k��g�G�"{d��>췏��$���z݃0j+�d�2�*�)��d��Vu����nu�3��I���u|!ؾ�C,G����4c���^��Wn��p�+��Ks�YXג��pѓ^p��j�`c�ki@�V�#���{�f"��fL��@M��U���"��O5a�&�[pH~�N�r�Ds���]��+<�,\2qy���u��캦�ݫ�*����Da�eI�	r��ޟ@�@����E9r��,��C�k���
8��Ga($��sFZm��9��%w��`�� ٣�-j�=����4{��G�	�=�2�m��t���m~k��=��Y���T���`'�w�4۬��n/V�sg:�Ǔ������cn��6?�W$Yv�0�{������^݂�ݥ�{�vU:�\>w:_lr��G ϰ6����gν�}�j�«�7Z+�l�3��]��c,�&MD"E�u����10zq�7�oJL@;�},�����!F�M؊�~����� ��O�$���F�5��P��*Ŧ��B�a1	�ry]v}��[�j�I�t�Q8�/��-9��f�$��d��Ϝ���GAhOO�԰����#�dh��nI�o.��q�VѲB��׎����>�N�U��:_Wv�Љ��#)G�2c|t���_�V�2���Հ����
��ݯ�:xrwB~W�+�>��IOT�괉��@��E�Z/���FT]Rݤ@}�i�x�H%}�Kv�i����FT�\-�s} C���=�ߜ?NV'Lqt�RE��+�@�/��������QG
������ԣ�`k�����?*y��	!m�wݭX����)��-�G�M�J�3���N�q��	�@�B����mµȋ[��,SD=���}��o[���z��XY��6�'�������y���� ���������K"`-�T�ʹ�\�kﬥ�m8��2,(!,z ��\M��n�������(���A��@c��������sWޟ��X��VӋ��#M6��w�V����c�!o�Յ@Cא��/�nB'������t�i���bg�m�C���ZWgq}�D�Wm�]l��ThI�X)��o�m��;&�vt9v��!��ށg���4��>y[�9�È�w���]�����G_�%����J�Z�2Go+)s��ߒGAHƻ�<�g�����Ǡ��2X\6��s�W`c�S���w��oZ��9��ݿupA	Q������3�5�5I� ���^;ZY%��z:��~5��L؃���W�~������^�I���H�J���j�.�t����D+�>��Wf��'a�9�� �7�|��qշ��n���Y���Zrg>��?�<o�*���-�c�@��}'�;�ˌ��F�70�Z��
�c\L�)h����)�`�ձBwk�Q9�#uSU�<5�WOrL�M��������6R8; �UBO�,�ܛ񃬽u���5s�sa���������o�,��)��/1[�7��I�Wϱ�k�Ʊ8�7{c5fI�=�H!fYi�u�<�Y��R�I��[-�T���2&���a��c�1k��w.�u@����m�)z�!}�>gI�%*TiS��pZ�x'���-���S:b�,��<6REB`��XP����.6%P+�򶈗y���zTv1��X�Uq��{C(Ԡ_����g�� #�vf�åL��<$ί�T��ͱ4 �5���q�g�Xo� �x?�d *汉;#�e��T������z�=Ke�Dp��Tқ�������a��\� h�TKg�bS��U�	_�W�N�
�G+�H�>O
k�e����������_}���4C���
��L[{D@N��U����U��]���Ҁ�� 0Mdy���7���ޟ�-�}7�/�)�qzV����(A�.����ۂ�m���`6/�V)ﯿ�f��?K:�� ���F�_�|��<>z�X��Sr:~�?s�������Q�癫��3��9�?�@)�bWU�;����Bu��~���x�����֮\��ָ}�L� o�OlKp<����)�@P�`'
�&�ïBr�Af7�[;�2X���|\f�ľ�lycS(F��o�O��q���4����2m��ڑ�2���%�� ���5eL�^谢�\�q�e�Q�8�Gv�����D���pѤm̈́�}�[އb�9Ȗ����%\eOZ)g�_�V-=]�C�sr*�q**�5�(~�ٜY�AW��Z*�;L�8�0;E�=�^��=�:�d ��,��W\�J8s.Nm��b���RH\@��`0���z����x/滖J��I��}�J�`��I$߭���[��4����A����1�B^��|_�գ M��}[��5���N��c��)�y�q��%���_p�j)�+L���GɱUtͮ��ou%j���Nw�'��DM�,�}	�%������s�Bڒ�?���k��`+XiBB��1\'RKz۰˔*��0Z%ܼ�D��n�TIG��~[��x�:vm�04mM|=bK�F�u��{�a�~<���,�Q�gV���P��{�V
c�53Pg���ӳ�F!�\�
�C���	�D��N�}q5�eO�6�^��n�Ɨ���%�ߔO���fn���R���������c~ Eܤ��i�j�k���m��,M�\.���g��(�V�r?��	�3����[���q����ى�!�6h���@��,;LZ��\y-4םn��	Ux��:��C5�2�4V70O���3��x�~�Cj�~
�����L{
2P^L�?z[�qO�Ƕ�gso�UA��������p�q8��h�w.R�����}�\Ƥ@nj~�G[��S^^��~��kX�~9Ϲ�C��=�`�ܽ+�Q T)���Sƣ�L�gud�N�3����p��1�(���0${��$��Q�0wL�w���3��Pg�X16
����Qlrul�����&���qt��k�(J��2t�s&{"��,
�?/�bt>b`��-6 ��L�T��pK���v�x�w��ƫ�^{n^w�_�ɼ������jWU��PJ2�_���x��p	Hg@ �\���*ފewD��wA.�Y����������1b��Y���r�mؠ�Q!�w���9!y�WR�]]�4���l5�k���.&��O3J��������zs��m�([�s¨��N]��]����b]wu�����.�A�����4m�h����Y�f9�>�]f����Y}��dR��ݜ�;�Ѭn읙>˙ܙ��5(�/�G���s.E��}�O�����`�쏞l7�u���=�m9M׿�;��g~3P���|:N��[`�Uy�` ��<�5F���˗�D���S:�������(R��38���&����:�(X�c�״�r���b�㨞��p��q���r�i�]�]W�6m��N.fg�_����e��wKCQ`��5+��I���Ӳ�_�4��F5S�� ;��|k�L�kɠ�$N����g+�_[Yw_���c����P��j���M�kx�a�.��?�&�4eg}�?�%�!/W@��;~7묞��.�{H���xgG=�����H�5�t��f����gIh<_ťH�p
�,��ǉ�l�ߺ�ZQ�W�W+��f�AP
$�GU4���������1LW����]@z�\�����Fc�Yо��m]�I�b�<B�ݣ�`C{��l�talc/W�k��r����ڣa�ȯ_��.�VA�o|�T�R��]+���^^���R.7����NGAF����0p����~O�**�p�6KP��bcZ��ľc�ݫ������&}�>��5%�&�NG�A��"/�o?�zSk�Y��,^��w	H�O2�pF���M�B\>�9�t�<��X����d���Q����6ܾ;� �I���{�;�s9�t�5�X13(I�򎳶3�W��I,���}$�Q-V�������n@0�~K=V�o�9��N��p���pO�����~Uie��έB�Ϫ�n��[5j4���
{�$�<���{/ ��}5�
�1�����}����ߘhFR���~���� "���]f���Oyzh��܁�����dA:f�&�8-�l��U�5+GW�Ŧn�ǔ�6c;�[z8���У��� V>$�,�!,ř$���p�H{,ǭ�
��Jߥ;�QקV:�ȮԎ$�G}��#Źy�MOgm/j� �fe���~��ڷu/\�QYI�f�0<ϗlҡ1pԧc.�\dCEe��`"�_�ٝ�?�ljm��U|l&�`�������_�O�
w)~�!K!>������{� �>��֡�O��ؑC~#y����:�7��Ɯ��x�˫�n�m��|b]l�j������0�p�u5f��$q�����c�?s5��aF���v��Q�ZEe�����qd�FM3�\�k�g��C�3

s7���8�y�0���N6���(|����y��\����߮�rR;����i���'0�P���k���;/0�n*�*�9�������Wf���X�\/N*�"3�Q`�n1ݽ��;{2��M�����u!5�w �������z��DKA2�￴�%�$.jf ��?TQ_Uh�>,;���a��8Lpx�_ӣp��]t��D����L�6�ߔ;,V�p[[|�;p3zx:���@:ciFf��2�A�V�i���{3�Dg��Bi�����Úx��]�Xo�?H���5h(c�d�A����RDTg���J��Ŵ�@�؁��ǰ�����˕��
M2V�|J���	�+��/,���*�N�%���fal��fv� Blg�UQDI�Ddh�Ν ��衽��iD�,@!ℊl��+1��c�j���k��꥽9s]CAy��&�ye��r�Xa��c���w��-��\����tR�n�.�F����[�j!y�=Y&�T�=v��|ZZm�z�[�� �!��^dŪK��sk�\�]�#m�Ƃ��O��3����WB6�/8�e"ft���b����s�h���1�R�<���W �h�Q�/~=܅q�s�oɜ����nڊ��9�k���c��Kv��m����n	$��xP��؛1�{W�][w5o�
���� L���"T�23b�w���٧��:pZB��K��XA�����rĖ�V��	�E%���lw{{ڽ ����^9�<A�����l��PX�=��LM,��6�X���Q�fh�G������#�����&�!t?���wu�� �6���~�C��7<�LA�m��:�5�逞�v53z`�ؽ"��=��{<G�p"��X��ę.�T��ml�[����t�|,�GM��=������0���l3��e��Kxӣk�RO�>/f�����Z޷!����T5�c� ��G���M���L�ԩ�H�q%$��2|+{��4�a�\S����	Tf���<�������~��ٖe
ד�6�^��Y���G�'
�� Go��r�0�}N)�LL=��n�S�f/V��F��SB�������Lx��~�h�uy��Cah_C�]Z�H�d�W9KhuϷЉO�D�\��0�k�jD{(]��6rif{/�Y�E����s���I�"������pg��P� �]��������V���O�	Z�%qUH����ĵa�t��H��?&����z��cg�r�������j��w5d����)���R��մ|�N>o�O*�d�f�0���ք�L��e�����#N��9e��zT���!8�8���˵����t���:ɶ�i5
+#�u�b	G3@G�>Og�V��u&�8�W�p$%Q�J�����e�& �0-�t�Ò���9��TgN���g�=��_:ʷ+��7O�󾦎{������&4�aV�m��<P<�'e��:.�Gw'5��D�P
6��l�^51����y�`$�kt�.QH!�-��_��6]O���"A�]g��KҜ];*�(dsT\�����9
72��`AÓ�R����p��\��B�蒳��7l�}�ąBh�U���-�~ؒ�Q�����&A��a���Re�����sJc�𞘒�'9�؆�p����ѕ�J�7��v
-,оH딏�J��݂�X�ݳ��uxTA�R��'��+<g�m��46���i)�x��y��g�:�P�\;����VR�m�����(����D{�j�N���	��¹|���F�l5�%��M��J!�)���مf��r�V���zQ���ܑU��	ZYk'�=*�ҫ9�(��08��d9��=�Ӛa�ҥf�Ik`]Q��S���"��G�=�ݲ^V�F1ft�y�<F����,e��Lo���ra\RN�8��ս��.Ύ�`'`�P�l\�(��(�]&�s��2��0��{��>�s�u��-��3���%?�����L���<���ë)Xx�G��K�� L�!��ӈ�C���*�Ůˍ(s��j:p�3'k��K}8q�����;�e2�	�L��x�.�����]QMj�-70�-]���o�T����m�n��d��
����4b��~�n¹.͘�0vή~�W="&|RЏ�(��O+2�M*ͮVjp*ld�qj�n =o�z�[�Ʒḅy�Q)��
���:8�@�l�X;U��aN`(�~W���'2-]�Ye���n�Y��#��;���M	��O�0���L��CX՞�Y�.o��P�a�uM�S^��3�Ԙ���+Ov͙���Q��Cw�NT�-z��Rh�8�8�b���3]go�E ��|���1�|��Z�����!�] ��)s�S�ʟ�_;5J�a���c�f�{{�+㼴�]�6�c�*���Fo�7Gő�#�����*�$������J��}��a�ڮS@�� ��_����?j�
�����(��+���8]g�o�Ʊ���Z�`�eN;C�uk8�7���G���\CDD�>�冀� ʻ��+�s�ei���۳�)��#��m������ �h9��W�_壞�YF�h �SC���W��8���[�ɩ��e�\�»ڛ��r���R��؝��$�(����&��U���- Ra�ȍs���ћ.��o�T]��t����/\��i?��A��Mο-?��n;����.Uȶr��jh+�s���X:p��W=�Rp�L�g���J���Y�e�1�ܹh;�8hi����q\?Z5�`Rwx��'�ws3=���|v`�К���n-�܃�)��|���un^�1��k�(|3�	���Ϝt��;{���^w���h�W5&�L�F�3�l5�kU�^��Hb�@ar?5n�뛚�����3�9 }7r�r�.�wt�%�GF8o���Mx�E�:ߌ��HRaI��R�C�Oy�x9� ����o	w�(6-����i���I�������eXK�6,8��%$�Kpw����N���Kp	�����ۻ�y����73��W��NwWu�-k��n��r=���W#�dXz,<>w��-+���-֚����а��8[��'v�����t�>�#0�}�� ���2m�����=�Au�'�g0ؒb�Q�cj�{k���kv����/�@�C9�geM�it?��+��6mA�>��G���R}�q֏_��������V>(���tśP+#�e��<xѽ��ePƶ���f�I�VK�c���9�!7��8��W�=P:�#�n����P&qߖu�\�����E��Á9+��wQ�q|xx�T~���hߑy���/7�'�@Q.���W�PAT�X��.r��)q'\Wp�B%r�����L�����]@E	�����h�w��m�|aP�gNM�1���sIx@@�uG��*otr r����B�l��A�$w�cژ��e�q#�&�����Gt8�s���I��j�J=������*#,������o;~p�m��yK�Eyԣ�6: @E�]5�J?:��r|�Eae���k��N�uҴU��� �?ƪz��"�n��u[��Sx2|�;A��i���DP��_Xh0Y%Ń��{1v��$�/t�$&����:�hX��;M��'���@�9 (�^Ñ'�a �jه��`2�"�_N�4>�)�%x�~I�e|�>>���C�SMJE�]2�Vc���a `��J�3��Y"f>`�lk�p�G-
ݻm�BX����I�D*�U��_/g���~(�ߵ:98$� ���g�Hg��d�h�F�L|���T:4��N���8~����ŧ���t��D=��@V�ը�ͅ�+�E��B?+U����K��*��؀�Ǜ+�5tI��eк�
|=�ÿ����:,��S�Z�D�m�Y�L���DX���:a˖�����Dn2a�C�L��!=y��(\�n�zR�\k�v��itG� E�� �	k�v6n�[v����Yq�l��1��zה���Y�#�F�}�2����˖YOq��&ג�;�����VtВ���:͊b1[�ʓC�=�����"�����/bү4h��[��j0��I���,�
$���lY{�AL�t��[PB9o7+G�a�mb1_��w���Y�F�5#��^AOW�C�R�i+���#T�sj����Qq"T�X�˞���P��3aꌺ�{����wI�`�4�'X:�`3�cqz��	��'O�
�n������Q�硭�c�/-�T��wbL�1���y[E	�K�v<�Lu����5iz�,)�Ŧ��O��� _ǯ��*v{��ȹy��
b�f��^K����>�W��C��k�"Ր�퐷YgE�4��{��A��L�ۄ�=4�ݫ�����Vr�k��`��gV���W���[��)���۱�HM�]J ��.�H�d$��6a���4��y��� y��}�I����˂hs6������ĥĄ�&	��̦�'G�v/7�Z���WfD��l{���>�}�}mҙߪ
E�`�w�� ��1�ߔ
���ʄc˓�/ 2�o�@������ˑl2yPFv�6��x��ɖ�A�hW��+�IUrԔ;_w�O��'�̀��lp�TU��6�ik8u��@���cy[l��9��#n0�M"�i�����~���7K��S�|秃N��{��:}Cg�Y^fz���DԦ�J��b[�2�KW�0���6�0�Sᣟ�-�M\�Zd�o��|�l����T�g��6�����.�N�o8^�.�{<ZyC��}�܊��5�~̘�2����Fx5vR��gR<uCmײ'sP=\��c7}���[CK���f���vI�c����W��-�� �!~����t�����G�R���a	(���=�]YT��[j	��\շnIw���ݺW�`�n�����ybU�(���h�HȪ�m&��<�ʹ�O��JϽ�_�~X���R�15�~�מ��=����c�O��D���FT�J�ex0QJ�`Ϫs��[�����{G�Y�eSX<{��u[1(q�1�t��z�d�|�ṳ���ږi;�Y��ב��߫���fý���2M�~j��܎OUyp�^IUW���D��g\��t���?��CDL���/�1[��K�ξ.�&:m��{BL~��7%��u�@X�nj����􍸛�*	fu�h0I�s�m�0�� tD��M�ۋi�G���];��Vz<�]O m[��Eհ���ۼ$�A?y�F�h����K�A~�!�)*'_�ҁ\��K�YPt]���71!,������4k��S��}�B�~t+U����˼il��C�j:_�ܠ���q�]G�U%�FVW�P�o�Q`��ـ�H�,B*xZfV���2S[]O�y<��2�x颟 �����~Z��Yw�p3��Z����ģ�+U�	̵�+�������vzj�ӥ�'����7�f�%b����-AV��t�2'�d�t�ɋF�:��YⲺQL�c0��:��uq$Z����˴��^L�K�
͠EU�m� ���Nӻ�:7�',�/�Z�ڴ9�g�9����c�K�-fh�Oǐ
�7��e����"��VL���C���(<y�sy;�be����-�09��K3K.�����l�F�d������"��U�j��m�V�][�^�����[��ݯ��6/�G��x�y	��Z5�T��B������@w���޸�V߹W���@7�%�k�8]�W�6h��Fi�^:WW�Թ�J"C ϙ�h�t��>XL�4Þ��6��ws�uw�n?п�?�q���iE_��$*�L<<�h�˲2�C�6x~�P7ف�.[�F�|-u=;;��-�+d�A�3B�2����^�V�j{�89k���Hv��:����of�[ߴb��/f$z�����,&�9�cġ	
]�5=��

¨/}�i�UƳ煭=pa�U��v��������,����?�wY{�t��h_|b��[�}־�$�PBUJ�F�������>���t�P��r:���}[~?��J�y�92�s���3���A�P!E�GX?g�|����DF��UG9̀��+�8BY4+����f������AW7l��Nv�J圫����p(�Ϥqy#�<�g\����]=Z��px�n?ߥ���5hI��lbWi��n� �̃6d���ބC�5P^���[��V����g#>	���z����d2ۮM�h�Z;@E@�__�lתҎ�G�&�@͎_�}��`V5����.�:D:fL�-=����;�����b�!$����?5IT���U'�=��oh/�5s��S��{���]�6�\��}��MGK�kX-r6D��/���3���B)^�Q3�|��/P(�i�xw����Q�E��1��y��ը%kgQ��[5ʙ�4�.K��_0�6�xP�'t���nG�R@����E��۞�W��.Ǻ~��P��E�2QkV��|�5_��r�"j	r>>�LY<�0�i���~EG�h��9I�oi^r�>�?�Ƚ���b
|j4�)�p����?�J����N�}rǁ+23R|�`��=
��q)������u��R���f/�ω�0��8P�S̎����܇���~=��<%ᨃ���w)M����ۘ\5�1��(s1E�����/��c,�|a���Zx��h�K�H/ s��[�V-���(J���7rH%b�c�}%�g�i����`��n'5}���H�ř3��@s̼�/F�wp#��h�Î����G�l	���&�Cj
_����/|��v��?|	�ì���?��g�H�,'��t��,�5�kŞ{�H��c���q]Ƴd�W}�x^q�B8��ᛉ�m5�Kf�X4��HZ�%�����m���[�R�8����z�R�z�)�R��v�(UP` T��.''���Rt�����]��,$��¢��������sJ��Bs`_^-/N�
��vȽk��K�"�u@�;w��b�ph�ۧ���Ok�>��3����V���QJ�ʮ\��9������D�'��YW����Z��X!��3�mS�����w3�4��N\���-�Mglm�ډ�8�{�L��'r�]3�}�$	���D�Eӝ����%���[ь�}������� ����e���@+ ��To������olȄ�a�d�/��%�bf+��z �͕�g���:��VA�X���cyYܻ�3����e������5~&�G�(T,�8|���ȅ�<�(���:���x4:q�J�g�+#���4��}�D¦�����:���B:��8]�oͥvt�Q�0��V������^qpF���N)�<dA��mioId�(?� �n�y��ː�u�\�>G�����ͣ�U�û�����_���ΛC�z�܄=��BNN�7��9���ež8ޞ������1.R���P���*&z��15�Ӎ\E�'�=zsPw��fB���Ug���P��b�xP����a��
�~��B,�n���M\�:�'�w����>�m���5��N  �Į��I�\�O�����a��Z������z�!Bl%��^h}xŔ��������(�W��ݢ�a;�T���I��u?��&���+M#�	ԩɹy�8���ݧ�Y�/�WT�۪�@��YF�S��T�߶���]Z�a�\�ܼ7��9��f�5$Į��� �/Do�5�{wc�_:�9�'J�i��vJ���)$���d�T����Ӆ�f+.�8&���]��>�u����TY�\�o�7Z�LImï����z&�pL�����Kk�t������{P]^%E�޿��m��f���w�o�[�Ѻ�:*�b�Y���"B"���0_�]47'܃Ѳ����r%��T��h#�vY�v�=�KE��'����@�.���L��o�� E�!����;������h���p�c�^����#ӯ�fg�f7g�A�xŌ�R�;�T�����7*�W�6��G�xo^6q�)-��{�@wۺ-4�*w����^�7�Ω�.k
��$�����>�(|�/���$�'&�m��â:�J5�#�� �_c�:Y#���:J"p���)�u�rZ�*n@�?����޼��h(+�}�F��EF��c���XihkX=��4t��?à5���4�nT!r Z=$rd��c�<�>		�o�����mO�#5:�{�|=��gJ2�.����%�o��o�����IsV=�B�~��<4�5��]f6���W���n��(���o�+`�Fs�@b��J���˂l�"����	o��]�G��k�[Oy���Ob!��f���4I��L���I4\�6-H���L�?�M�2� ��]5sk�p��f�ݦ�Gb��� �LX��ĭ*o����]���]YwS'_��M�c���޲�F
��k� pFK�r�/$Z�[�];Y�gV:Ou���@q1a hϵ&�ÍI*k�*)�0��YGO�Uj5����6+^�س������r�+�����b��O�|�{#��L3���bX,�'��3y��j+�oh%�3�?��0�� ύ�N(E�8��
5���wz4���,��,�����s�$q���=�3���=w�@0�Р�]����=��j��RLqjaO�s�x��t��=������٧�Ks����eO,19{�A����a"��#hх�s�>��������iyn�K��-�pN�]�T�RG���= \?��C�}���0͊�<T^�G��4U��t�{嫇��_�"���)*��񅙇V���"+��>ee�fy�&�Z,oYh���i!wN��F;3[�W�D7��ʹ�a�Є��`I��{��2�'��D�o��W��'WoA�̊�R7��C�/L��A(+��夆�/goZ����p�����K0��CXb�_+�g�-��,PH$Hr ��Y{�L!#�X�\���m���7��<R�l�Fn�F�T>/Z'�N�M� �b�KHHL&�#`\�����i�=�O����@�	{*�?�C��<���M}(ğw:T*?c�m�%���_���)R�g_���;0Ռ��4�T2���W�|G`�[[t���(@A��Λ�����s���@��a����l��N��a��8��8<Q��i��E|�,!=dԏ����xj�&u�2��A�	�����۫�yz,ߙ��p�8%46oD�r�RS$
�h�����F�"���ƾ5�{���z�����N{��M�*\��j����@�
UdK���hS(��?�������w���Cx/�現��)�������Ј�&*6JUr���8׮�/��):�Y�����W5W�|d���G9��G�-��q,��Ti��q�r�[��vJ������,�Hhx�<{l˘r7��6;Q؏2�FX�P��~���RseP�u������JAhp�q��_)�2Ę��$���FqtY������`2K��o��%����-�rv�7���Ί�ф�3턉���ᢠ̛�%hŤ
)�9�����I�0��!���ԃ);���㖤&2�5kv��w?�r�c�q�}!���6-Դ�؞�:[��>��N�GE���w>k�{Ey\+����'�-��`�X�1˵�`�p|rXQ�4bn��[q� ���O\�t��z_�T��F�=gu]�N2�D�܌����x.Cz��.@�R�v���8��w�J�ʋ�7iQ�~3��PN�8>>�"����YmԱ��:<<���U�n�1<ě���|A��$���*&���(v�<`��	;��=��E�۩�0�{����[��\^%�xC"8�+���~w�Ȣ��׊���f
��N� ���c�6�I�'�_�����SC
����Y�3�q�IӦ���i���>,�P1���+�1�4}���7��4NԸ�Łؗ�8CbE6U��(d0jcG�i`�թ�\��0��A�<M���0��;�]��1�W?�5:a�nx��\��+���qT؀@�(��tPj�dk�t���xF�ĵ�����.�^��煩�GE�;ez�о�}�u]Ӽ�����IR��ϑ����ײ�7�)ɣ�6]�^8Mj�+ɓ���J���,�#�:t�Ap;��vT{���~�ʢ�ݽ���z���_��~p;Q
��*�7�4d���'s`�-l��'<��*�������R�
��ح��;k�՝���\�F� �/S��m�ll �iD�M�h��B��!T��8��U��W�Jg�h:�u���t����,��@琣V1��j���׫w�Js�ph���>���f��{��o|���y~��&Y�F��lmkk�yϼ����d�x��)�������i�m�Tdld3�!醌%���t��g�;��B�H!�����,��7���)���]k�����B��Nh��Yϯ����|�`,�5���q�Ύ�u>�[=���o�Fw䢨��1�g�����E1�W�+n@�M���0�	��f<T�U��������N���^Z�3�
�?p���k{�=��UIv���3���b���|Y�^�q{�(cE�C�^ ���z���E		x�5�V(�^Q;�J��������x���������&�%��eb�|�_���/x����kԛl��W�l������1l�E"���rG8�d�w�~K�L���:��u�]6�%cҨ�A��}�Phf�-ZnCd�sx�O�U?Z��:��c}$r|ܿ�V_#��q9xCuR8E���"�7H�j���lE��S�퐩��騼� �%�]��!:�X���X�˔��І�����'>Eb�8|�Al'�Ā���ԑ�j�_�2)�S��^Q�f���>��v}�!	pF�paQr96��m���V�Rg��x�x:���b��;�_��7ԙ�\+��,)�+��~_�`۫�"���dWH�qPu�Ο�4��(3[��K5\�/gt�������̮j�wRM0H��nO9 Imt��[�Wԋ
SPZ�]�t�6��H�>�n�%_ ���������-w��/�~�1�>�YI���ǬTK���ʫߤsW�Lq�j�x�l>�@d6�C=�E�5�~�8�`,LO�G%h�}�g�(ˣ��Y����{�s�p	�����l��}�a��B}��샥�9�-����_���4�L�?(����	\4�P�f��/��e�V�O���f�Es��-;���d5�@���tPmk��~�˵�:�c�6&�q����o�E{m�Z�=q3��0�`�rL�]A�^_����#�0Xo�D�fj@C�Zl'�H�^�
��u� l�e��S�h�[>cӴ�Ԉ�b�B���@�bCx���z�0��\�mmMf!��<	#�?�a�D���P���)��R-ri?���3����
�H�~�B{����H86��{C�D zڴ�fu������-��5�	�_�a�+����c��t�9�h"uzvk��	܊pn��V3N�j��9�2A����j�E����	�WY��SqP�����A\�����^���N
GI,^�'|�tOpokx[՝�[���ٰ�#�.`&���q��J�,�(�,r��+��<��Q�A���ݑ\tS�Q�^r���B���z���M�U����
���`��Q��1�i�o�ZY�AQ��賰�亇UQ�[���1l���F�r�Dpz���އϯ��D�gl9�a�b��o�M�Nm.�{:�8P�ۋ��%��w�hmn�)*I�œ�⮆��5��n(�Ј �L�u<�����:C^3U��]�$�=8�7�����ߢ����ΧP=�8��wo�N��a�?k�hs�z�u��@W���^�r[|��HLpJ�yr����s�5N{�3N����n$Q�_Ą8PCɡ {�n��a��҆p��B�I(�%���PP�܄��Á�����q�L�3,��$���8�5���!��v�bѫ�R��%c�.�;_��/�;3�҉�iU�t?���:;DyJ7�ƌ?��t/�eP�*��6��������6*e'�e��G�>~���DP}B���E��y��vE���"�O� ���Yw?�����"�i�Hz�1 c^�<i�ߩ��8qp��U/7o9T��H��A7(�o&>u�R�>H���kf�TC<,�	{�]����=+!��,?">�m�`'�T�j��w���e|]����0_�������'�,y9O6�ƌ����˧/2g�5"��oߓ�~c���rQ����/���=
]3^ҁ�`����?�II�0.�VzLw\Fl�'!)N2x�o��)y����+<8Z�퓘�T�۰��m�X�J=~Vpq��W�������,�s���;�٣ߤQ1��E�C��Ҙ髉��Ѯ�m�"F|+��B7�,�tq��;^?�O��{�~�� 1@�ai�(���"��s�^�qŪ2� e���mS�,�'�g�T�������Ng���� ���cԖ`�ۑ ;��Y��u{�[š���9�SA��#���;�[r>w!�p+
� �{��x��-騴����-�~'+EW���|��_�}:N쩁n��M3���W��9��]0c��;�������-"���&f�f�`�8O,����P�O��	2��B&eg������c^$�$L��?�n7��P9�v�Ѽ�$^ ���B��T+�@j�����Z����C<����O�(��^@���>5�a�~�Vd��6P8_�CR�q���4~۴%,9�ء�*hkF��NqHٞcT\{j����<mX��?"9߾EɚΡW�VU�s����9ڄ��k�v��T��T�9{���	.h���}^�k�wv�m�Y�g�r����bNZ�<�0�bl�(�;;{�s�	1���f�E�C�]�:#��PHv*�~�=0����j)�+J+�P�U^��@ğ���Je�߻�͟�"��c�H�H��1}��y=8muI�r�����Sj�K[�1�N�ٴHR�E�-�t7ݳˬg锑I�G@��$= ��o�qsV��g�������&�؟���}�v[�%�*P�'�myO&wX��}�uH�F���X����w�Ӝb �tB��J��5:�]�J뼰��hH4�$��퇰�Z4�~K-_��N��������O�{��PIk����"��ʧ�]���dH����_����[~p<��ϳA���i���v��Ѿd�9�-�y��L^��z��q��d��A����6����he2֞~�����$��J�����Zb���!oЈ���f:��9�`x����H)�-�A�hF~?��m���2zt�'��4����N�M�p���|..i����f[e�@Ց�Զ`���7����(�)��J'�]z>��L�'��M9t�C��9:N��a�����;��\��zH:��%m�h�r�n=�Ϧ�>"�L���LΫ���;�pߴ>+n��L,T�4n��H"��aA�L9S-\C�����*�vp����/^�
�ˉD#����AizA�
���B�C��F���4�%��H��������M_x�}d0V�NG}KK{�a�|�0�O:sdHB"z�0�]4���;������EF�ґo!�%Q2��2��7�q�ժ��"���Pl��C��
��B���-`�aW{�\i�bg�q��s��kG�^�$܀mY�.`�Wn0��P��n�~�:��w���i�!��;�PO�����5`WK
c2����馩�ܢ�P7 �a����םL8�9�>�g=��w���?v�L����=������^|s]#8��m)*?�kk��n�]�,�� �9*���7<�UǍ�Qg��aŽ��o:=�RƦe �t�\ɲ�Ʉ��7-w#\�|#M\�[ ��g��c��|	����b�# ��~}�9���<��J���k �/�z{yX�h��
�2B�p�`��?��y��0�&iz� �8�c��4�(sVH��4Vpެ
�X�x�6`����,��+��������}�z�� � ��uF���� a�G���!�.�h��x��oz݁k5����5j�Т��ھ���&R�>>������Z1T���D>Q�,���b²V���^�������ɵ���p�Y���<
��˜J��&L���G�E���MqG~ge���C9�oZ�F8�V��3��#K�g��������#S��v.y{�/y�5���	��<Ll˦`5oi��c�����bf����\,�/㏵"�2���{�����iZ�:�X'�p��nd��@ҕ�J�m���u����[d0rث�EÝ��"����j��h�΄�������I���@��:w��$�T�0l	q���OV$�SW�_���T_�(��|\�'��H�������{3�v�c%y�x�SN̥�����y�oe����ʩ�;<W@�(
�l�Zkб{ǜWev�4����Ԣ[���������IR"�>���P|���J�Lv�{����%�K��������۸�<y��+���P�B�ud�}��μ"x�5}�ѠT��T��&{�W->���UK��(,X�h���kI'�d�!��1�8<-h+�J��jU	��zY֛.=�+0����@�Bx})>[�ͣ��Jo�����B�zߐM�3�D���сfa���]
+��<��SkQ����:��U��>�6�l��-�\8���~e�i;��#�<F����.o6R��>b*��"b���Z&�vCh�qD��H��d�R_�3G?��_fLW�u�#1�yx_0b�Z!/������o������9@C�,CAJ��`��$�5��e�R�=�7����gM��E���s�|]�;4�t��t����Q!���u6{!%�/���ܹ,����{,�ע�/=�JQ\�B����C�Ih?���$Z���=�QoR��d� A54=��]K���ZE&T�� ð7��5���e��Ɔ_�Q� x�^fC�B*醶:�a; E�ͮ��*�2���lgJ@�]�~�G�>�����e����TPi��V�9L3�&s?	-�ś�� e����qR��\��m��W,�a�X� ֪9����Pӧh��Aw"1-�1K.|�u�8�>��V�H%��,��kbe\��
~fў�	���O�;���I:$T]�[��<���uq��;�"��R���K��%���Z��`�:�b'fR���)a�]�4���A�D9w=K26�R�{y؋�MC�?�M�ᕿ�����}���y�>��h:a��_����t�ބ��[�u:�Zy�'�#\l��Їy�����Z���hG3t{�O;�Q��t)���4C)�S�����������d���)��J��|�[��@�|�5_�i���<��q�Ky,�؄Hou�fP}G�2��Փ��s=�lCz�ߟZ�k����2w>'m1T�cۉs�s�Ň2�Ǫr�V�K�*���1s���-\��y�<~z�g�a���U�;��������4��a������ic�ܮ>�P͝le�%v�{���>�P���6�r�hD��{q��n�U~���	@�:P�|�3P4����]���3MY���<���|]��cI�����0ts���58 p�g<AJ�"P�?OzKf�fKRf��;~:\���e{�9�_M�ϟev\r�ݏ�Q��Z[���uĝ��g;+輻���H>��{\�2��	]�w�|F��Q�ŵ{����7� ���f�pЬ_��֧O�Y'9m7�]��m���f���r��`���in�ϳ�Jb~s ��V�
NI ���+�4t��]�>��v��$��p�{>��|p���{;9�h�\� m�;�;�ha�w/��c�6t������E�z2��hɯ�Gx9��=\� � ��V�NnQXmj�ɖ�[�
��c����
�����oU:���_��ڮr9��� �E����B���U��)8�t��0��k�""I	W˧4�<�Y�/m��O8,�|-pLJЍ`�7�X�q���N?/{gQ�����,�C��4P [%@l���	�9cu�;_��%!iސI4�ǀM��Aޡ�g��c1��O3%��$�S�8"���c�����i�\'��{e1E�+j ee���?�Q�]�k��s&窈3����6^�L�ǧr��Б2A\�S�6���k�Ŀq��RG:&~�L���S!�ѩ��͝H�L��_�
@C��8&���Z;8��,�8ӏ�D*Ĉ:d�-y}�i�;	p�Y����i�9qLS�~N�L/�=��1���PBMW�sv����F�l�F�j��ʤ���2=�Ѻ���ޮa�M�o(N2$e{�e3�%���
��#�{7�4-�}��["�Ug�\�g�W������(j�Y|w�}q��'*� ����:{�G��$�MFw:Y	&��%������2#������S�5��9~	P�% <��a��H$ʸf(��W��E�p\-���R��Y��`�e��G^�Z�N����YqQ�w�h�/  w�u��8�>��z���݉�T�����;�ڟG�޿�a��g�-P�������M��o>B0�wգ�W��~,��}N{�&i(�Vp�� ho׾fN�T7Z�0�O2]Єu�ٻ/�U72Qh���Jq5�؅��;Jl�(�����e�� S�B�������+>��X��֟'Q��H�H�t�O�O%���!�@�� |_4���L�Ƭ�\%�Ň����`�x]H�RY��(�fo'Q��W9N˩��E���F ��� �|Zr{�ܰ��VG���Ɛv�\!�6S�k�Ѕ���	Vw�ӑ��J��Gћ�L�j:^%d�B�jh8���G��r���a�՜��Tc[
]��\A��+��\�m=e$�SWtM�Ƣӵp�{�\��d�|�,�l�1я�cQ7���hd*��}\("�\[���0&���>����b���n8$��h�}�R���%"����GI�9'�p�wb��t+�w����]���IVO���TLo��eRz�2%�om`Ŀ*3���L��,��+�h8=
�VZ���o�`��|�-R�+�/���� ���s��N~�x�8]�w=�d_V��V�B��/����c6�Ys��v����0����
�`��
r�m:|�M_�[�-�X���T���+���I���\�ί?���V^�i+jэ8����u:0�Auc��1�ty�X �p ���U�jz8�x�b�Pu9�жu���Ԕ���єi�;[y9�,R(ƴ���P_�v|%0l�C6Ou��ih/' �͜7-�B�C��}Jo�����$��(��(Թ������x[`%�q��a4����y$2�I4�(�͚�]L~T�	���+u~����_i�N��X���.8�t8Nv�rӮ����V����D��%�G談�B��/i-�Q�m��n�N1�G����^5P3� ��3��`���z��g��!�$nE��k@�h��?�:\E����Ԫ��ǉ+f[��[��3Yl��m��M���/�낳����*�4B�LuJZ�qm�`Qo�t
Z�*I�z�l�C�S��{��C7�Cqx��t�a�&* ��>���v��	�csc!ć���s���D�������<�r�W�Y��,\ơ6տ��@In�?Ԅx>7v�B�U�~�{	������*T��S�~7���i��4�"�:K��}��N��|]x��+2�D���B�u�n9�[��󓖬���3���Ӛ+���V��a��x���6(�9IT��
��0�x5�P=�r�
��yb\�ҞK���as�t8��+���i%�?�:���R`8iѶ��'p	��B��;��
u���d��+f�!��u��Ҷ�NX@��3��5_�ް��R���li�/�M�@�����2*
N#ۢ���-	���'|e�ҷ#���[�K�m�^Ü��"��F�Ճ�]���uؕM
�����Fd�E�u���}�3�����>���`;BҜS��V]�}Ft�:���zd��	;�2�X����`����;�O��_����(�*&�b��e���`04�z�kƹ���{dnXz9ag��Z���	����h��k^�� ���]x�Ľon�E3K�ל���6��f�?���J %9�PH2C�<���y�G����\���k�t�芨��D�E%����^�2�#�8�I)�4�p7n�'V���7��B~�2�#���D��S��t~m��l5:�;�7k��L�4��k���wp����?�_��>��)qQɺ�;��+�b��&i�R��e.f;�%o��(I>|��Hks^��Lj�!H��0G���T��7��>k��dD$�ܚ���/�a�'?-uQ��V�q7�]tn�t\�hO����`\y4� �Ԕ� ��(���-�Z/�79�b��Fή*�\¯���=Z�����y�ѥ�"�5�T���d��Y	���g3�M8����-�n=�Q;w]�����f��7S�N��v�yi�����m��5hk�
����2Pu�,h��@V�qk����;$�5E�l�쫿 b�[ƾ�LG&P�~�2�C�Чs��C�:|�x�a���{�^����};(�� ��Xe��Q\a���H}=�f6<����&��]�(�&��T�n�J���撆R�W,�R˾m� �m�f���8\H�lP<&�J���^�E�hf)�>jt7*�a:�ԭ��w�_�_\��G�n�%�>y�.�*�=2��2
ڵ���v�'�[EK��i"��c�V�4�^�v�����߮$���y�"�U�9ĉ>!�����tVq�}c��0
��m�A���v���BU@>��<�5Q�N�ya����w�]P["g��c�ͯ�q�b��D�y�jSk����;�+����ߺ��QutCo9*yH_�U��UMn����mn��J��"��/H���S���Eo�l���0jh�9
>�gb��)��Y��|̄ku�pe��/:a��<F�
��g�~Ӟ�$@�(aX]���,{�_0B�������>N���$tR���҂��5[��i��C8\	��<�^�r�s�a�r?|�^��f����nⵐ�M� ���M�F'T�&�d�A+{2
^ן�t�<��S�u��>2s�2��+�\�������l;�w(��$_����}} =XR^�7nk�A��7��ᝃu�m+���LL��Fg�K��B�&zk\�+����|���Ptx�*ԛ��e��Vo��m�8�Z܁�f.�:�朴�?@)�*,_�9b�������\1w�cW1l���`t����fn�=�Q	��Z�c��7��ʫ^O��^�9���I
6Cn���-x��C��(��W�\D#?ꂤO�v}���'�ݜ���!yj�x�&�G��Z��&����黊����]���L>�gܨ1�2�
v#oj�!O�V�U��q�sh"���/(\�7�ڭ'E#b�HI�"�ŕ�T�F�s�x6�Y%������%n�┹p�K�'f���}��@
s������O�+����+��6
�屉Q�Ŏo���a�0�|�\e��6V����ף�����M��ڦf��}N��5.@��;��#3���&Gk���K}Ul7�����t'u)�P�4�M�g�B�W�VA�o.S�%`K��{��.6���a\0|ƾ�n˵!�]L+[��fpǣ@(�j�m��::9�Ԯb�V��}xUx�.�A. N�����u�E��9���UZ�{�6v��:!r�R���{��C��U��J�b��<'��Aiz��[�(�}�Y-VC��N�?����;�J���Ĳ?BFq� ���u�B���i��/~��d^��&`�Y�Z[�K��^ ��Q�v�q��T'[S+�Oo�(wÖɓٷ<Ŋi�e�ͩ��)N� ��"��'ۛ�Q;y���kW��b�-�Ŀ�pp��ާ�G��¥S������v){���eT`�5� � �% ��� ��w��[����Bpwi��h�����~�ٙ��6��z��[ϭ*���g�	C���:	?QV/�Q,In�.��ϵ�.�����͵ͼ�p%^�L��A�p�S�PŘB���焽�E�o��W���p�8G���Z�eRx-�J�UC���}�
l��3k���d�����M�:����)
�?�Ұ&C}�WKR����~۹��r�0n�W� �\؂��nzG�cx�aid&C%�'v[�2�\ei�$2�0�A]��;E�[���!b^��n^�0��aP����Gކ�h/�����6a���(�E*�K�Fl�b=N�z�y���&I��W���v����G/C�H���&�8҂dd�� jk�h��hJ��;�E�4��w�Q���I"G��Ƞ��û�6��z	� �:2�C�� ���k�E��A���lݾ�/�|���nK�Q(�:��%�ټB�,&���L�J8��>�?� *RPpXJ<��sG~4��:�Yb��ᙧ����.�*뎎M��$�<,���|8�u(�>s��`?��<d���r�&Rm<��W%�?�>*��}b)�G4�S��\e6��g�{�O���-+]咤�.����������c�Y�=�����S̯���,Lw�8f�T~J9T�{��׊L�s��ë�_(��zE�1�iD�1����T֐��\3i�%��o�CIA�G�E]no�����h����:��� 2���[w?�����5������]1wha|2�'v����r��k��q6�/w�{R��a�f-C4��'��$a(V��-�1�ܹl��E>�AN*������.Q�f��U�U����	%9��2�AG�7�11Q�s��W�˚.O�f���>	o�� �y�~��A}���7E�Vy2mŵB���Z��ۢ�58�1	3`+��Y�����𴩓*s�[���y��2�lRB<��ʅ�B7����iuϫ�������OG͵b�|�T(8R�_cz]�=�2�8�K�g �Qӊ��0�4��k�<6$���`!n�U�$H��{���{�b��3��b��Q��T"���%�B��j$�� �Nj�F��C4�� 4��A�.�f˛n���d�|{G*��sO�A�-Έ��Y�)rx�k��P��>L|�+P.~�!�>�*u�*Z�������.?r�[(q����.�H�k�	3c��`R�ۜĶ�7���מC:�ޑ�B	ܶs�א�R�u�!5	v�(�O(q�%1ypې
(����Dv P�L�qJ���=�hq�y�5c%;�V���I��W�B��&Ƥ��q�c^5�`��n"vZ=d�~�Rf���ߘr܅�k��%_a�+7�����$.����c�ȩx��|�Ρ�g��u�Kn�-駔)���QK+�s��yñy,��Q��G�K;��qO��v|R8r�	>Q^���V9CxZ$6�K7�!���/�����Q��	��Q��z��X;'c���OG��h������kY���!C�u���e���~"�x/��^C�Q!~��1�A�#fK�D0���+�k�*.��jT�rpT��4�BS��v��%�m�J��3�f���KT,�)���j	�q=�1��6�=rLjD�P:18�!ysdKפ"��R�*�fjT�TG��*��2[x�ʞSv5��yߛ��,IU�~"9��,B@���d� Ŭ!�k����k|�2��x��,��wХ�O{�3��G) �^�`k���\��`ȿB�:�6�)s��� 4)� %[�·��d\���j猃�q�J�>MEƲ2�ɫ��'"��f
K�o����J���u�0��N�.�x�Z�o�rm��M.�Pu-���L���������v]2¡ޚ��o /o7(5�6D2�px�#ױX�e�M����`m��~wp>D�O3�� Ш�ZӔ�p�S2���m�qJ�ڕ���5��5��_���f��ґI^�%�N7ۓ{�ߐT��!S <m�N�[!I��\��q�R���2a����@n��i���B�s�B�|3斔�o|K��`=˅%��>�>��U�6��ߟ�H�l�h�V�n|�F�X�:�v�<j��aj�
�Ʊ@iv��i['�ޮ�13E������,t�]��JG��N�f��)Ĭ�i����>�ʟ7���:N������:"'�s��R�����J0%��%w���S��"�����B�8)���Fq`���K�-?�ܫ�{Ӿ���D�	�\>EK���@&L۝�\-�y�I�}��m5�<q:�F,.�/�W�Yh�Qަ�����ǀR[�^g�x
��"�v�k��d�?�~aR��&�����c۸X�i�@���2!��k�C9-g�F`������]�ĺ�S�?m��U�9�k�I����P�	�o�MjNU��>�$�v�l���ߖ�/4Aϯ䩲z������,�֖�(���P��d�%�Xg��/&���H��UlP�[:�Y!�
����?���~E��fl�78��cΔjҏ�H� �h���QL�.TF��a]� ��w?M�J�*�>h����<�ߋ����I-z�I�'� ^d+�z��]�1�
^X�h�+Ť�������!�� �	�8g��K����Z9���fm��F���(
ޣ.�^����k��7��O*T�C�"�-;�W���@�E1����ƺ��c ���۠���q�MF�S�>���C5�m���F;������M�!�˵�����s`��/0�v�]�z�D���0m���L���*|CW�k��Q�b�8�x|�r~y�[���zht�vˀs�ީѬ���x�����%$��_�p���T)!D:F飞
�(�!�b`�$<v�?�i��{��x�(�\`?zÚ:1��}�X�{�}���!
�( +:�,�{答5��0��f���w������
�BC�	,�s��𩪷T4��S�;��"� � �"3Ϥ&��&JU�+T��HV[��9z�^��^�On�q���V��;���
��MF�0��`�R�z�(�?����E|B4��n���u�kv��I ��R�ǒ�ʞ������t�.��|�X�r���`�<��7'��u�o��/^�P�	��H�燝v=�/ͨ�7���@��ܦ��� i#.����(B�J���m+����N�B͎��(�b�1tW���1<��Z�0��Ow���:f^#��,+V���L�P�7�-�7�M��w�Ü����c��Bu}��.'uU�߷�����GW�����V�E�
1I�5��d�tAFe3��aYIY��*_��a��2�I����5�Yn
�V"'<L:��f<�*�f}<�8��)�KvXI�E���\#8�c���zg;T(D,�s�Ϯ�8g%n(r�0&�z��W���fd��B�I��S� ��-��KL.�W7 +T�R�q(N+Q��ˣp�<�]��J�ɼ�£�͊{���R�ψ��O��8��yk:�hc:_�X�1^'8��h�%T�`y�y�h(�ң��B���\O�}_𒬪�/)�爇���P߮yW���/��ss|�?�;�C�,]���ӧ��.+Q֓����xĬvO�É
�U��_I����j���e�mt�;e�7 ����QY�����U��������U����r�D=�����l�s.s��Sϣg��FE�/6&��IW����͑w�J�+H�m�V��)R�"v�u���.����U���oxd������y���ne�:\�:�5%KՏP䷸�D��B�wP4�)[O���r�W�:´ā�e�^�|�o�h�-c��D����/L�G���b���3�ޙ�V�4�9��_Two9c`��t3�_�4�uR�Mm�{�1uZܢ���n~����'t��z�2g�|T��d��:	"M)���km�����ch�֮�#��|���(��b���ʘ��r�XSI}�z��}�R�k5Vl��^x5�I|ܺ�pY�>�*�ެ'���h�2]H(��#���m�#�>���.�<���7�]}lxb�+s_x��́��
O���9k�D~����-��F�
�����ڣ��V��$�F��F����v���C#p������L�M5MwM�;)�F��-Nl#�<�Iǉ(l�k��u�_�0߼D죊8����VO�j/�Dhsk��J�S�R�g����K*�&�A�؛7�F��n��Z�+�6j�?�O���l|�!�-�[�H��6�NmR��\n�R�'|]o�UVB��6&�0=((Ĝ4�(��4�c�>ky�-����ꉽ�Q:�z�_�ݼo�y[??1���ima�f����'��z��RD���+�F��W��p3_V�H��_�8��f��wj"���<[�]�V�p���/���y9ρ�=���aC�F��<�s�Z���������7>�#K0b�T��t��`�,��l��{���W���f��"b_��F���W� �8Y�$5����.Qǘ�-�4�D���Yuܾf��D.�d�:۳��8]��z��k;�z�JR����y��HTH���kT��譁��	�<i�e8�o�&Ϲ�¬��Pg�?�O���1�>p�}���+�|�����hy#���ǭ�~prt��)�j��2�B�Gz�pM8��s� V.�El#9He�(��嬳��&�ó!��&Tz'S�"�[�-3��6qh[ZL�V��NN�_���89]���1������ȝhv~zzw�
�2E�:�Vt9��Ӛo���Wp�X�+V׼��L�v%Ҍ���c^T������V�=��U�ˤ�`�ޱT&R��_��}{�P�+c�r��*W7+�(�08��q��wxS6E-����Ĵ�8z���]zB��X�qJ�aL�d�A���	I����B>��j �����}���Uvi����St�����Z$G(B�i3�J����;�:���:�����Py�0��U���hg��5#���ӓ�(f"/��L����ftO����WoS�4�������*��-�(�έ笞����J�h�,�"Xg�7>Ӽb�]%pUu��Yt&b�쁆�u���:_��*F���Gy-���&VK �c�uA������Љ�AA�����?��'E�
���쀫��:Zԩ����b�ߚ,�ĳ(��oe>n<��yؔ>�}���RKh��%�/��m2��m>�G1�^@�
Q��>8���ļm�x*i@�"5aJ_���t�[���E�w���P�Tfr*�?������J��z�!��1"����qqyP|��D��cmZ�D�K<��wUy��"�`
� �=�r��B�P��Ԥl0f���*��2u����X�wX��}>h�U\&�1rݬ���G5w�~A����G�����>���N�҅���*l%Ł.�N�j�lE��:�
�|�պ����ٴ�����1_ac&�v���[;_�H�V�m��� 뼒A^U���pflf���Dv�h��:��o0�����xQt�h{��2�#�~��S��9c�?�-[n�X���b��\�EiW�`��1� ֢b}��l�s�&����G1�!����o����������Ɩ�6g�*�A�����v�����6��,�����o�}�]T��P48��u[$�%�>G>j��
�gD�$@�����s��o�(�P��em�J�Xo|5Rǣ9�_bG�c���3.2ϯ?�X�?�G�oȜ؞�{t�&7��l��\c����%M	�J{.R�[5��r������M�S�����mF��ͩ�x���q�v=����Z�kƮ�
7�u�*�����kg}o�ְ���!r��pPё��Z3��t������D����fMG*��ڞR)<��<�ۄ�勰ᝁ/`�T.Ұ)�[#&̠�V��C����h�l%�I��%�>#�/r�tj��NS�J�/�N�2W>u:ݽ!	u������cmj2�q�_���HvL쭈��ȯ��1����z+k���
:c�	pQ�8���C�X���c�����bBl^3��.`���,��>!f$��E�r"�ESFqQ8/A��9沜�M�)�FP�g~'%g����p��s��R	h<B���i�?=]�)�L�#��I�z4pvn�z��YX�� ��x���?I�\׵���.��6n� �
f�I��t��U��y�[F�k>��=�}~K��dxe��8���ם��_��7�n������8P���"K/4OTJ�11�������/�F��2M=,cj>$}��IY���s�sVW�I��V���QQ1 �q�!�/��ʔ?ښ0�~��m\m�r�t]�X	��j�i��y���S��k�4�p^��)��Yz�1z��iXF�Qo�c�������o��_�ot�۟:8���+c`XM�����/��Fl-��ak����o[�#���9�ߟ|��TC&����6�Lų����/ÀM}�ȑc����S��	\G\��-�M�I'*�==���'��
9����5������1�QOxN������/TF�̾�����̆�)�S�d��+Pb�����4���}�Mx�*���n�V�25"xH� ��m�y��WZ�By�h�	�G�l��w��Px�։�����s܉���
.?	�3�Q�J��Ʒ��J� H����=�2Q�����E�����җz��`޴Y�VG����Cө	y���Si�@��K�Ts0�Ķˤ�u���@�	Oj������7���8/2k7p��R.L��a3`H���F����6Q�I��:w��>�� ��$~�)��e(8#�8�7�/��������5L�O�5�0��ޜN�#s����S�놢8����?�'2�v�k�.YF��%��6M�h��2Wk=d��+��za���X<K$�\�+j>sv�����W����S���۩�b)������4���mk5��困�&=��
�y_��7\%�N���Ǳ|�X�
�k�
�T�r��#6W7S{��XP�"��<����ղ��}���Zr(7�K�>`:i�:�2�5�Ps�h�,��F�G�9`CO^�b\�3d���}���jt+j]�l�;�|�՞3m���+����:��	bLH� �g���sS�(�)W�.2x ���g��Oz0F����=��J�||��ч�a�q�=×�?��U��s�U���c'AP�.���4��Q�a�H�U59g9����\9���O�>�������mqGTG?~,�7���l���_�>�r���M.�ծ����?T���}�V2���X��v���K�M����TY6�7/��LJ���E�5��H<�\�D���E�7?k�"2�dDpG�^�2�t�+��\�m�aݺ�kgI�\z�����>خ2����և1��]:T���p]��_�rI�F��=5�Mőf+e=���\��C�e��&��ݭ4ٯ�Қ�߿���;����rU>93�[����V,����wJ苄q�o.�.6b�8�k�Z.Ё	���'r��8E��Z���e�V[W[��RD[�GG$��''��u3��=X�j�`���83����#���~��*�U�ԭ�� ܲ�����	��{��OB箣�3�kh�e�f��� �Y���������Yb+����n�N��Fݱz�A���@4��t�����r��z����g`phQ��L�#��+Ἔe*��3���^!�Z�W~���%x�4r�h�
f�F;�slQ�@�%�_D:r�m%֍�.��?�O:����۵3>�B)�5�O�ZAX�s=�����'\�"�K�pZ�ڟ =,Ui}��Ӵ����~�]��p݀���x[����f%I�x<�R�~
�t/�h\���i�8�d�s�K�����u`L�0� B�7i� _�D�u�C��J�o�� n�K��ޗN$m;��D���fZVh6�hrV�i����4DS�\�&���ʂ2W�GjBCB2ت�H^"�7�9a����2fr����������DAz��UI�|x�1�e��p>[�nܗw�~��
�����ΥϛO�]�V'䒽sRF�}�Ҵ�+KV�V����͆K):����/�O��W����ޝ�=S�Xc�K�s�u��-��s>�[�G�C������/����V�j�n(�}��kK&���LL�o#Ԅ�>��P�:ll�RKR>94�d�֌��'L�N�f�ƺ����TRQtK�l~�⪽7�l'�׊y��NDm4���h�t��&%�1LZ�SҾ���m2Gy���3(Vn)�5O�������3�I��q�����b����Ij���D�~�j�g'��4������� �T�rN��=" NJ�ing3��²�:@�]S��:/0(к�Y��z�aFk
̆�� ���i���}��hZ���`�����=׆���(���"�j��Q0��7o\���16!��������Y`�����Ko��r��j!̥s�����M��8�`��7�u�@�p���T�CWq�}'�`���^�L7

�[؄���<��ԎT�P&n��i��=j�|�M�����*�R�yT��k����cU���0%b��R�s��I�rK��������(+��⽯N�K�^��7�G��sAB���Ӕ(��Ae����8#H�������� e[!��Cm<�Ӯ��s�����'���3�<�8�i�Yʅ�?������o`�z�д��JOi��|�V�Uq|qI�VqS)/��mӓ���g�Wa�Ln Q���Hᩛ�~W������ �����/�-��a�~���yv����p�e���uB�p��]"]��>�B<���]���ݐ;)��ش]i�%ߩ�����2!U�&��ku�&m�.q��a7s��9h M���3�m3��k�a�?��b�>�ŋG
p*Q�v5�v��fM�@�şܓpX�\���<�A�&h^3��81�|Py� E�zhS�˻<���&!t��E�h	�U����P�=��	v/�c�{�1,���O���Q�����&��{�v��:P���>����&��ѓ�s�$/ў�P�K��J,.���ui��s]76Z�@īH4�xո�Ԣ�	qx@	
	1�/�j�`��� � P������~�mH%Mm�\?�1T�!����^��W3��^���""�{e��1���͵s~cs�_mw��,z����H��矒�^+�C�r
5�������6)A�g�!XJ݈/���Q~�~�S�@�y�]3W�d�*�����P;B�c��}�l�]���;�(��\��l���i0U)E	��f����7��Y���V[�Wk���JF��we�7�������zU�zC.�`����P<r=��M�<�r�f�{68)[�/����>���~�}ڹ:-��Yb`���3�ު)+Qf��$ч�q�iU7+�b��'���G>K�)R6����א�}+�y'���V{%)��	ŋ���Dd#9���x�?�]���t������4�}�?�:=��[w�s޼�U�.�k�|�"��8y����"km�l�7U�դ.I.i�yj��l�fj_�7�+��|���9���<��.�oBg���Փr�{&��$���ր�����h�H
2����>Kv3���Z�i�Wς�4�&^&��"�E��\i*��04ĝ����Sd�C�d0�]︧<
w���4�����u��g~���:��n *<��)s^��
,sP�tS��2�ǻ�Q�V|�=*�5�8���x��c�L�l�ٓ0Q�թlj��W�޶|��Ϧ�[�-���4�5;A*b��x;"o����)=��5?�����*�~\��Z�߀�;��w=1=|w��76 ;�`D�<
��v�F�g=�%Wo2!�}�N��RF��JwZ�9~� M�)z��7jo�X��k�}°�l]WPy�d�e#`Z��JF�0ۤ�{����jg8��Uń!0���f��?�hɲLS�p�lu���k|=�9tL����ڻ}m�=��>W�7���3a���ҵA`�CQ�il*OS��Y�D>�]ɞ�|�0�����Q<oބb�q���PQP~7X-���ܰw���iT�/�e�D=N�%�~Hc��(.^D�a�,ޫY)*�*��m�N�b�^����C�8��[?Q��-%CusUK-��}��mi���rs\k9G�"���9KHo�b�~ܰ`��'��q���F(���rC����}���Y['��mNH����/{�ޯ���S�-9/]G]K��2t�W�iw����9J�ŵ�ǆ���I����a�h>4�݂w%�h�{0��d/��r5���Hv� �3�1�!� �/�wM��
��<���iP��ǝ��n�������X�^�:Mك���c,�~��ථ���f��U1�2Nx�,�zU��,8������j��`50\������\}����<�ȁZw'��.�^{GOvM��3�E?�W�;�+\�uҧ�̲�[�&�rZ|��Nc���u�4e�j7�,O6�Q�~䤜��yu���y��<+W��Z�2��E���uY���D3�61��]b�>�K��;\V�����Q�{RP�B-�S1�!&�������9s�w���[K������}���s�U�q�Ps�R�L�5ok�m�ti���k����q)�h>�w�n:~;}�� �����I�~����5++��)NN�������m!��O.v��˼T�'���J��-�7�&��(?���J�eQу�~�j���ڛ��ƫs�� �Z�H�;.�I#�)��q�h+P�GEC�C���9�'����^c�u�Z���Mb%	�]���(}hbz���)��6�h�׵t��[<XB��MB�X 9l*;�Yҗ�g��t+��k"��Ч�����#H,п���3��T�Rm����L�e
�@�i�'|���K��������U?�F��͞~W[�X��Z�>��O%"��k "�6)�˙.y��}c^+�S,ɒ1�@̮��L��(�:��[�>ܵ�'�Z��U�ez�i:��xF�u�˗����.f'���M
������'���5�g�2
��+�U!��bm�T5+S^'�+�.�v���?��	�%�ݾ+�\,�jc_ɤ�������/�jM��ZUwGS(U�|��?'���ǹ_�]�D
r����{	��"��v<���?Cv]�\����҉�%�O��=�z�Z���{2� �t�37���ǒ6M�����l:���M� X[.�"�A��<=��$R��9|%U�h��d��)��UFA5�n�j2#�q�O�����~"	1N���y��vx�5��Uұn�gh�6~��6*B:��Ք�Q��V&o���/-��It֧w�k2�pi�Z�敉��5[�_5������&�s7^>�����z� �Q$(�E�q����%��S��E�i�y<7�"��oS�С⛼�����������]��{w���OwkU}��E���k$��&-�h#�~���⽩�ÿ�>���z�d����c;�vq?�&��s����5F��ꆐ��k�����J=zᇳ��t^j�ts���)l���r���i\C�ސ��ܗ��/䴅{�KX���,��ڼ�6RM�s3
�/Es���R�1�@tC�WYI܎�Z��P0����W*���ʭ��Z_�G�:t7zպذoUM�.ת��p525�M�Z�뻁&q��)���ɪiO�}������ZO?�G��L�A����?��0�e�?kr�Ԟ��'L�H�,�S��
 �gHG$�-�;����o��_+�h�{�{G����|-~���6R>dv;�-��8eZ�<_'�8�Gc��P��w7 -����;����~2���P�5�"��o��c���J�O�,]��U>;��[�8 (���s�2j���t;ܐ�%�2��ӧ� -�0/�-�^'#��ϥ]h��t%+�|ؐ���S_�T1�u>��]��q�F�W���G"����c7��N[pX�ۯh�(K�(ɯ�0����Ά��GD��u������>� �g�zP~��z,��â�c1S8��~i|w�SJ�����-�B%^M����L�G�Ľ��i�W���s�%��X�?s�	[�4��j&N����u*�vj,ܹe�@��<��qi�2��^|H`�X��gll28��_��1�$�PjJ&Dr<��G	M�eν`�6n�$~!F�̻��2"�(�w@��[7�}7�-�o��8hg��2�Q?:pl	vh\!x�Җ���6��}���QF���p���0�>v�k~G͑o�r&����}eve	n4�!��S8�����?��[{v �`H�E�D�4z��ދ?�i�k������c��ht�f���\��L�S7ƿ����q�[�Xiؕ}���zhq�o~h�H,;W�ML�f�ѯ�E�ʉg�/9,��ؓ��6
���]�]�6#�#!�M����࢈�%���ݸ��� �+-��Ӝ6B˽��f`�6@�&�f}�� ��ﯕ���;���6׶�AE��9�@�w���3D<<�����䰀�FF��AA��������i��@44��b��d��� ���\��,���,�$p�U��Uk�����J��T ���5�͞�G��DW�����}�-'�[��
!HR�ն�����tr��;�/3y���q
��fg�GQN�{r�gh|�Q���d�y��'}�7��k�$�i���T�����H�Z�̂�0�����m8�~�F:�̈́A�)����NU⋮S�*Ϥ����*4���o}�¥�;�
Y�'kr[Qq��T�񣺕�:��+OI����m���[H�����>]�L6Ef��3�����1K�Ԛ��e�b���:�����Iv�p��9�9�Dteg��l�R	<�4�
^�ݠ� �[�����y�ڨ��1Y��:|�}: s�<�9�͈�xW
/n�6 ���#,�eM�� �;�� ��jX&�f�D�E=�/��!�U�����8��]	�7B�w똾k��Z�ț,|�7�"�7��#z||�����-B-  ��Th9W�	噾��P:���,��9���?Ǚ)��w�����EL��b7Y�����]L��������H}{a܍]S&�f��}ul��o�Z[�<6�����F)X2�'Q(Lw��Q�M�Iq�B;U6M����C:��-R�0���3`�I�v@ҍ�4U�V�؍�h)�q���qW�mc��r�zK^�WQ��o��L��t�To�Q�w2rr�C[E�;�Y3LB�eQ�ɶOw(�4]x�-�}j�3�B-�ڱ��g�/���+��U�t���{��Vb/��Pa�jkp~�������!i���%��kA��d�D"wBGc��{�d�)a��^x�[�\�g!���s���@<��͖þ��U�EN}�;�R__�@g�>�._J���P{2(w{|nNBl7���&��Lw�t�M�i���ɡK�-�Pz��:p5���q��Q��0;�ݢ�Z�S7�Rvړ5ǒ�S�pk�ھ�II�+�9p5#�g�C�����z)��^z&�W:��r�-'W�%'$�"�BJ����TBB�����G�TTT�<���␦fcck�}��H���~`��/���P��m}6y���4dtd[_>5]�E[��y��C>���ID�w��Q��3��	����C�-R[����\S��Є�+�Å��L&��I�]��X�n��Cg�J3�=����G�h�b��0��S�l+x��~���0� �Ɏ[�	L�dn �Cxs�_���\���c�>�>��e'Չ��ш:��s��e��'۾�L���@4x:������dS�K��@
%D��k�����B��
����[�偖x7]�h���#�#�	�]�K'�S�����Q���)V
TQJ���B��5l���Ɠ(n?>�G����Jϴ���7Q��C#���-R����q۳�x�L~X�Z�<�r�蝑�Ї�t��s��vW�4��s�M_�=� ��W�ʶ�&F�oh�� Ym;�#'���ȫ*���<�:荭�j�As��I��������唿��ӑ��^fQ����9#�<�L*�j]���Q��6�MqX�$"��l"qg$i$�QG�ה�M�+M��d�^��\��4��<J�(�"]i������A���a��Z7I4�]�'+l7��o�N���z��?�4��*���g�.f�������b������}g�˿���.�m���㘵�_�P�����Ⱨa���JrSi�n��A��j�q���EC�jH݊M��I��n�� 5��_
�|Z� B��OC.3'E��c]6�N��?��Y %��ʊ�ﮍ���%�h��_̍u����I�\?]����z�n���Ҫ;'�otM�H+JpuiQ�6�ׂ{��K-�j0��Z-ؤu����,��j�҂��:��y&	��|�d�}�
%KnnyDe��"��Y��y\�B�j�Ɉ:pK&(�HR�Z��n���T�����sr/�/���2�H�h�����@+=B1P-͙���NE����fS�Fǖ1�>z�/�e9��.}!�;�$�@��'�8S�5�XF�UҼ�?�m��}�֮(���p�35�n�� R8)U-~?�^��t{��'��a���f���I�葳�ϼ��j|;�D��4C��65���Wά�6/��� n���h��V=�߈��M����"����jڤ�õ��#�?н0hgV��I���2hjo�Ѥ�5�dI��0��y��KiM�,w77QV�<��E�iL��zI�9���A��5�±�K��!��jϮ���l�9sk{CC�8xp�q�֫��}�D�H9�ާ��j�,3�[���sˍp!���,>�Ą	,�m�f���\�iŴ�Ԩ�ܕ�n���l��tNi6��u�z¸v��< ǫ�PL�z�%|��3V�u?�P���v�k�ܗ�9N�����a�D[ӳν��/i�	�Q^�C�K��(�{k�	�h���E���-��5f�k���r��ə,g�h΅I�9�[u�a�ޫ��$�WF��� 0�ڷ"���u}�)D�����t�xw�h�bc��Q~
e�DDR4cV��Fk¦\�3�v���"PK�uC�Ƕ�c�u�}����5����)ӣw��B}g�b4)Y��W��Yt�����,cK�W�yp���](t���>t�ٶ�MV���r�W�h�^P�~�T<� �W����N2�ML��k��!�x�J����G�����׿��'>Q=�<���h��(���
7�^�7Co�X�F~b��:ڃRs8wzH1K�u�k�K�m��� w����>��ݡ����X��#�䋥k��&?}�c'��2���W��ɿ^���wO`Y1��\��Y��,��֞����˧S��*U�<0(�x�r{�V�|�%-���m7660	,V �KL0�p��^ױ�������1P���;J�a�4[n$-�����C�P.�SB�t�:%Om����9��W�b8�O D�R�����A������ظ�'���ʱ#1�5v�"QD��O؝����(��`��B|�&b=� ��M�-~�"�
X�_Ҫ�z��R�ɖ�v�k�#��P�sT�"����S}Ev�auN���043���s��ϧ��`X��!��?�K�bygƐ�h�+��>0q���*�Q�����Ow�`�UGu)$��	����͖�2A�S1"��RMÍy������r���lQ.�߇�4���������b��<�j>�We{�+��N�xs
��u��i�SY�Y525�J��e6�{V��hp�(<�<�a���eQ�n�s�3H��i�։PD@3Ț�/����9T!�����;��.e)�J��R͈���$'�O��_Y�J9��8C��1Z�(Ɩ�*Ǘh�p��Ѳ�%S��X䣶?ɀ+>��l%�)p?s��%��f�;�0Mg{�K#�/0dM zu�8n���(�h���>.(�6�t� �>�oblu�tw�U-|'Fa,޳�����+SYI�0IH
Q#�veG���a�И���Bڛ;d���ڈ"�7=���̭���(�b)bi�3�쬊ǜ��ړv춄�54H|���9|e҈O����#~�tϬ���rS0<�gY�s��,�Ey2���E���u9����c�u��>ZTM�j��^}F L���
����M�Ok�'PT�+�f�kk��@4��ժ��ZJw�0;Z�_��?x��-Y�8$q�ڟ�Z,��ZRu�W�|����Oe�\�f�>��ȼ�ͦB6��[�X&��@�h���ܺ3�_��x�#Hq۽��v�-&Y��4��5a���B��iM�Y�w�	��p{���x�� p8�e���s��w���Cj�c���F���aT���j��lY�Z�����T���j��-8zH�b��N�j�f�J��>��n����O|�\"�(U����ǭ~uBcGz%n�c6��o��A����h�i�Z=G_���p���yИ[�My�m�g����ݙ{B���G���ȥ-#�!��/��iMONG>5�~}T-�z<�����-�81xx2Q,r�p�b��塄X:m%���t[秧��А�	�Sh.Yp���VD�b_B֐����x���-�`�����*���G�nARR�NQ����ݩ�tw*ݒ��N�wog�����y���s�9��k}b�u�N�݅��U:?�q�<<p��~�@�|oo�]��RX�\~�r��ŗ/_l��4�hx�+�o}���[rˢ��]��8��lb��Wg��ڬ���@�>�Y&�)4o|�z��8M0���y��M��� P͟1���z�њ����0����_胳�2Oa���|�ȗ~���=o�R�5���N#��k����n(�_�7��r�|/����{���,@j�8ݭ�8��]�ݠ�ճ~񩲻���$�]�` "�ׅ�L��):9��b��We�]�?2��*���ړk/aC��*\v9��/Pj7�����>~&��H��31����.��yS� ��������a'>��#�����&��|��P�cyW�^� MO��X�?�����'�{AP�83���z�8����S_#�އ���``���H-�5�d���俿�D�-A8��r"N'�R7bf��9�|w�:���G�441��&λ���K �,""�.��Z��W�X��l �)7W�����_����=�3�*>G�+˄@y��mm�-���짶��u���^"P����Ю�U��%7����`�j�I K��	�!��!�⸢I�&
L��"�~��U����MN�7w��T���S��s��,*)y�A(��A��ro�i�}��{ֈ{��ZJT�M�j�Ɉ"�8��c���7�������^ؖ�%^Lv���@���^�@T�5>&9�L�sVW�2��c"uť����F �0���y��Z��&����Vzb�`q����цb��&��|
�M�`@�!�U�ra�� wg�<z���$q�)'��~�3S�?�H��n��Q2���u�2{�n�����]m�撂�K6���}���Ve�
������͖��u�����j����)���|��^Bq�m�}֤�J����$���-.*)��U����m4�BԦ��C>�:�B����U<JJ�kX����O���Ѱ�t�:^
�}����3�9��4����(riq?�����n��܎��y���8I;�� t*|3����ue�x�-�Q��@hy�k�7�4���yi�۲����T6d@@�ͪ�)wT���2��"@2U5Li�,��|��#@Qdq#: �(�X�*�>YUxh2�|ȼf��EH��r�8��0����4?S��[��=���p/5.�K�}1���v�~O����(彮./6\�s�,'U�?���,ֺ��3ʷ��L&͊�ڲw�b�)T�7i��e�LZO�
������s�� �s����.tjv������'�dˬ��ʯ�D.C�]����<V������B��9�9Ȳ��{�;å|}��4�X��vµ;�f��Bj��
��A�ecs��E�0��״S�2���^>jג�oA&�k�|B��C,▎&�KO��n�Pyƾ�]�<��{���Þ��>����Gv���I�[��\���$�񜣭_���?����)l����R*�]N�]�Хް��&`^��q�h�.�%����a�Y�=��<M'�X�{K;�]	V�la��<=��a��3r�9��@�q�0P̈́{w�mϽ�6�F�ޟ���]���l�W�8�k��Mg=���Eo�8��?9 �d�Lj��qA4"�":9��|�ݤ�r������o]��jY}򔝼�U�s�;���u��x�3C��D�]nlQ�U����J�J;�&$�x��}����F�w���I�������^ ��M����m�� ���o�*�T��+�F�n�N�Z�:x�]%�o��ܶ#v\3}�,�z�A�Q�l�{(̙�	��s����	)u�Q�8�s�ڨ�J'ؖ5�}l�.;����ܠ<�%����v��P�:�y�yA�>mk:��a���$�q�=����U�~[�6ǴB"�o�ce_�$�4m[`x�u-�G������5a��`�Mf�goq�����h&6��A�f�Ps!ޯ�@(Eh���򺦍�]Y�"�B9�aҗ��ĳ�ʀY\��v ��J�7n�a��*��W@�o,-�e�v� Mta�K&lv�RY�/�Z��^�1	�
c"IS�,G�tt9SI ��;y�;�˵%;�n��g��ѩ����>�D�$�t�y(��BKF���9Uw�]N������IL�/��{&����Ɩ{�[��EY���7.�M�g�5d��S���?��]������
���2��N�-��B�����FW0O[R����]H����*��.�c�i�{�J7w�c�,��eY*��q�3H�U�0w�
4k0m�P	wX+����f�}��v�����S��������᷇p?>��^����l5&�E�v���ngץ��n��f�{�z<�X��#e�iʘц�4}.�w���f���\O:S�j�jG���]t��"���+��DiC#j�m�'L$A��C�8������b���V4�IJE����uM
�3A�<��$�D.3���hD⑿f6���7��YG��5���ë��#mmri2HON?[k#<�g-��qA�x���Khն�l�d�v��XG�~�'�3<~�75��{/S/c���9��y��R}��"�,�˽�O_?����C��#���(��J�W�<6Icd�R[�٫!J�Nᄻ�h��7�G�pP����D�����#�O(�!������#�}i���Ѩum�2��e%pG[��W��=�U�l�\ۅ��p��2��������F��G\��w�js���ڥd㿑��,$Q���F�b��\����s�nмY�fe��^Ty,o5��VRޓ}�o�)�1�f,���G���(��U�\@s�w4�5�04z�3>��z]�g�Y֝�ʿ����v�Y><<�I���&<<|:A/CXXX��	I�T�-mmJ.!o�FS��} [��-4Y��o^��C+�|t{(�*U��&sM�;�A5��ͦ���A��룋�����e~s_�c*� ��0�6�EFR����e��qK���YZ����$��J~�� 9H�_u�gھ�A�>0���A�O	]�^�;X�G�[������M4v��WFE^��_##��lccv���J;�p���
��nIU�{�(T�_��1��m��޺{���'W�V��܇��3S|�k���ux(�z'��X䩎��n�g%}[.�;��z�a�U6�?SO��е�皴�M8�C��.I���o��ـT�{&�$��o�Y5�*j\}���|��>����:�h8y �
��":�����%gs8���3�!�����~���R
��f�ff�ܺ紂��#?x�Po[�Ȏa\�M`�#/;ݷ���4�VG�`9D^ʇ���3�\uJD�,��g�&7�O�D���y���lN�������R�`���Xd��Ҟj�k�jJT�^5a3�Np�58��ǝ-*�g��1���+;��gP�
RdK%&_H�����H��_"�����)ۄ�h3�� �±
*�ٱ23331�i��:�Y�B3�����/}�[�-�l:�{��9w�xSh�n8������IáΙ�d�$qJ��0rp�L�xYÕ\1�������^jhUV�L6�cKY����ؠ����\�mVm���4c�k��l�-��\�*2�5b
p�ςZ�,��^�HD���z��h_��錘����I���U�YAܚ��UØ�&w���38)cŴ]���?lJ=Q�Q�$
�k�R�	Mw4MDb"���!o����j�:y ��B�**�b��d�l����Gl�+��7�8x���猷��<�Q^�Y� ��.#��ɿ�����ز�󥧆za��� �Te�CJ�[�r��Ǡ2�`(�1�Ԛ �F�6E�Q�-���.6�6IҦUt
���J̹u���q���
f��U}Oa@�2e��CAJ��0v�O�sC&�ƽ{�� �aȅI�Oš�0Ԋ��K>�^�p`~�5G���=)b�M"%r�=�R������3�owRп}̔H��*���#�3v�ˣ�	yY�S�N%����$�7�L�V��k*�U.�^'ǽⷿ�[������ږϑ �|�˳�Pd����m � J밭t%�|v�R�!$B5B%#`K���YZ_9Y?���^�������{<���v���-�GSW�F��`���=��r)+9=k���j��g	�
&�С�B����"�YӞ���z�A�����5(�K��ժn~���|���>�z2O2+1zRgVǫ5�J��`�[4�l���[�K���\��޸� =��V$!#�b�X�@��������ˀG�ND��O����z���PtMT����c��}�Kp#���,�h~�$�Q�;8|a���R�F��J���5���<��ۛŴ��J�9ayt����ׅ��ʎ����u���U���P�~ 1�a����J�ܩ����2����׀���x)8W��4f���V_����1<��p�^:ڀ��$-���u��f�ћrH��u98�S��Z�Cd4�R�K��o��Ku���i��H�a�����_�.�������� $z�Ԥq=1F䏙�&�[*�#���|/��q����:z�aN_7-<���+�����e_�Y?�_YQ�����E�"�è��t^�\����������F5�卩gg��˲Gڔ߮��3�Zv:�f:�>��ȱ�CV� ���{i�՟ #�힖d�Χ�R���}DE���?�:�~#)q_'5a�HJŹ2��*m��|�j$����V��oN����Z���o~/��kt��(Fݾ��Z'Nj��II4�Lש��Ǥ»À���^<=�����ҿ�E(�d+�X��y��[�y�{RqT'��L"xnxp�tt�&��l:Z��J-��j�[��G ��Ĩ��Sڟ���F�*��L�B��Ҹ� �����������J���W�ǌR��y7�#"G�_��DG��G����8��y{��np6��\��"&�m�Z�zr�8�@n����Xn9w�������Jms��1P��4�e�i0?Zv��]�P���B�7�a�d榪-?M�	m������ai"�" #�#Ee+���޻7��}�p��N�X��v��M�Kf_ճ�!�Mg���G�������݈S�Y�&f�L��uX-w��쭝r��F��r��W$�R�TF^+k��K���%�"�Wg��C��00
�|�����A6��@�4Zi�&}���rp�������%�j���mϳ��^u��[΋���:"ƒ+���:���m��?Շ��'[*Y�;<W�������Ar�NZ[C���ŵK����1zw�(�.�4��]�C����6�.6��{���oJ�;�f8�tM�LCEF��X����:�6���d0,,W���d�ʯ�Ң������~zj����i)|?���!<��U�;C�t\hh(�U�'�V��g�S��n�4��wk�����������U�s�6������[�8,���l��{"P8�f*CF����_w�x&DD�'t��lҫ4�V�$c2M֍���+rG�^ŕJ�B{����l�9.ތA�S�"�w/Y&���v�pb!��k����Ô�����>�]��*�,�N^\p�˴��Υ+�8?.��N��y+��J�z��;ֻ��c�
�C�4n��јݹ�LR��
�6�F�ʅ�aN_3^!�*ژ}T�z44����c����=��>��ȥ%-V��"��a��5����uf�|"L��<~h���
9K��{Z��c���kWW�1�&�+ ��N��}�W�����;�@�8���Ue�����z�FtU�34ū&�����#���j��Dܕ.��b��KA����"�-7��+Ҩ_���&ҙg���j���TN��ګ=�z�U�_5ݍ��s��h�`��{�!��F�b�dـ����m�&��Z5���0�>Zͅd����+l���al�L��&_����꽟Hf�@�iN�r�ʂ�̷��PK�}Z�w�,e�ځ�N�`����Ȳ|>�5���n����(xx��J��^==�O�=5���~�0Ý>l��h��!��VR�/nmk��?���i���iâ|[n ���pk�Ć=�2��QB�o�j\�*��jDK2	�S�2/��˵`��	*�\��B�de�ۀ��B��a.+�$��ot�P��TYOa��vl��t��Ά%���0��z2y�DH��('(/̄t�=J�T�z~�^{�Ѻ�Q��Lyz����N��n|5���+�������8�JۚiC^�s'�,��E|[�{?�
<�a���E*�Li�IW����.q'75v1�hV��K�R��ot��f�쌌ȴd=��r�ADd<$$$M����|��'�OH�"#1DDE�j2�l�FCG'cg�4!����ދ噅����gj��l���_�hUvGQ��y ��[j��am��=�=���uAi_�X�w�LO@��+Ă=\�t�X�SAi��ԭ�9��q�%o�$^�n�j��ƅ�'/M��Ȁ�wR;o�a����8�8���C{�u1�XeK;�P�!p�$Y�2����b,�i�4HՍWm�qI����ǜY� �iͮ;�e^e�_���ty��8�!cc0G�
̘*�v6��P#�T3��f��Ib{?�sЫ��4�ċ�޲��81Jݮ��w�4 j��Y�6���5�=�.?
]�|�
�M����aF�`��K�����~00�yJN�����S���8F���p��I�ܰa_W��)Ԏ����v�]%R��\��������+�[6�p07�$>Y0#Dܚ��Z�Rq�V:��:��^h~��$mNR�[���
�YM'��w��F��s�0���w}��VGg�^¤/�.��tw�<�~t^�����y��6��Bs�H������N�m%��h�:t����ʕӁ�FWsS�u�+��dɬ�8@xYV��5}�-$v��|cexy�8��;��&�	@_1_�۽�?�s:�����w������q���������9߶\�.\W�VK5�[�R}d���¡d�'�E^�.O��0U���)�=�w��ʹ�L� \.""���t���t�ǈ�vGOO�sRkK�Ҹ{�M�ׯ�^�&���wُyyy��-�����\�����Ёc
�:��$ �T`h�Ĕ7(�ѷru��>d���/��!�֧��F\"4Z[�ꡱA�!�0���S�qs'_u�,�s^+Q��.�(�W$
�#�#�9��,��۽6L�A��%?o��ȣ�@�e����q��&LH���`�.�僪BF���r0����@U�kĵ�����|�wM����xE���	W	k���[��+ױ}��d-��F�5����3�܁�E�'��_;A�4r`��!]���M�qY���Y�C�=�US6Y9�h�e��ec`��x��?���2�<fe�/���uؐ/��t�8.�����64*J�q�!�G�J����WLK+�M�k�����" �ix�V�~D%�����<&��38�>S��Ap��fo}C1s�
���C�p���+-֫6m;��~�:����}^bpC��mU��F�,f<�|�(
��kb1y�T�T������묷�݉ۖ?C�/2`�D��Q��^q�%��D*�C��#wx�7��K�K���$F�޻&��K�,�>�	@Ç"(��G҃� �Ν;��H�,e��X@�~�7Wnh���ፆ��u��k���������Ҽ�̴L��}-��H�;]}��a�<��}@���:Ar�s s�O&�"�^�Rro�e75���FDܯ�m���A�m�l�b����z��Qr;�(¡�?������C��V����1�di:A��B��N�_��]�O�o�'۩^�3g�����Oc:1<2�ZZ������Kګ{I&�fPU���y]����S9�r���8���! Rf�GZ!��.S[�~���E���x��q���[ XZ�.,	w�����P)x@�SX�W��
�13Ā�<����KUZ&7����5.�]�[G;�1Gp�:ty��Fm��A_1-���aҌ�Y&G��8�ck�a���+��4��z
���O&�_�8n�J2�;ߋ,��#��}�W���h�	������Q�!naq��JǕ[G�֗b�+?��>r�8�n%<h�!����$����*�ߟA5�FX�Vxx8 I_���նJ����(��̞�o�����]*�f��h�v�]*wL��Ȧ�Ad���x��ŕ^��}x���� ?R�`��ۂ7����w75�:�9m_�.��4D��h��279��!�9�r��Y�}m6�60�	�T�dA�b��dC�(oT�FJc�=�֬���R����̪a�~���|M�a�` �˷O�uK�+��^4ᔞ�L����ƅ��,��q	~�C+O.1.N߫���]LE%Q/5��Ay�IA����%�� BQLA!VOO�<��i�ֹ��*,�� �#�G�oZ�k#������={��7�Z��H��;�I�'��j���7[2�G�����[��)���������;�(Vm�
�`|�qbz�01l��=w�#��.���O���?p9*L��\��I�r.�ks�܍O5[dH����y$=��, X��U��m��i��z��ہ̣�+3�D�YUO��>�c1ҳ}�����վ&�lx��D|^\\\�E��
wh�YH3n��g0�s������;� �/�O� IM ��-����o&�� SL��:a�Q�p�)=JAz��a�	���tEG,�4��.�7%�#��a��g����S��8���l�,� �2\xx.�9!��:���`��߬#+�XZ���P�J��M�ˊ�.��A������
���e89�~49���RY�^(��ѷ�����Օ�]ʞ`����/����WK�zΓ�Z=K������ʘhXXFM��̊��Ԕ��H�'+��j�MP0��H�,bx~��˹ �d�|h����*)����l'&�*)@�	��}�3�����,>�m�졊�tF����j?����n�>"�yUjY�����Dc����Y�7Y�YJdϖ� ��pH���PI�����K��H݊'h�Wꦬ�}�w��12K�:t��k����:Ld��︕V���	C���I�t��Ә�v&�d���{R�+}�������i�D��X�A�xV ������b��$����X�f�1�sp�a���J���f�v����Mg���ɜm&�l�+�O))��;q�À@%ڣǹ]����F�`�I]��H#I�����k⣘E�������B�+����謆�فoa`B�*�IY/��r'�Y	k�h�ӓn��g�j�h=�_�y��CEȨ��S��,�A��ۼ�V�奏�����+"��;�8�>����ݝ�@�(��3:ŸK�ɥ{>t�_�wmpw��ֵ�I����Ɇ	����y���J\�g~�\����+EA����i'��n�G��t���@/e��Wo�j^��������E�����԰�Ild).�ف8�|�̌�0e8��ذ]��ӳ='_U�������n��Y@n�wmU��^*�����	V@��粧!W�r�W�qk���V.��q����5*8k$<`<���� j{5⳯T���T��b	����&��D����'!�J�
H>�{t�!�Ï��`�"e����67<,�tv�Rn�K���$f�Ea�j�����r]��`���y�����|,���;�W*�*�֡U)�/Tu}m�h3���H˵&���� ��pn-<>�����G{�):6��0ٳg�>��(<s7����ƕ�Ϭ7n��T䊋���H���~��,oUq>	"(�6|�S����7�I�nΪKܕT2'S��Id��ջ�K̛��7�e�o���^�7(f�i�],�0����k�Qq�����0�/�/��==Y��ZmH���'��W� �|FGk?0������撲�- �)��U�:s�zy���%^�vx��Qh,�)>+w�s��h�0��{�	�5���͛76콝�a����_P���$5h !.f�
8�қ@��y
�}�~�QR��6["D9�ۋ%�~>q�Y�;�#��`צ��e���F�Œ��s��z�e��]�2BRc���|�|��(��v^�� ���K��������j�U�ü���8� ܿE�p`��A�S�'G���l���31;�'�wr�2�8&VM|3���&(����
�8 ci�hhz�����b�eddL>�T[���������z�1���EUH��+�0*��&oOÛ"�9�s�����R�K/1�exR�87����2i2H��!�Q�������bnj�Y)BX2:͜%K�`�9�N��ɒ��@���B�ZӘ�FW&��Q�������?I	awM����H��⑔�b�7��L�-�bպ3�L{��WG"6ڭ4�tm$+P04E��	&<��h��,`C����� ����G"�7���T�+P�~�����b��ܥ$�w�XW��շ�͂vd���y/�1=\9�I�͝e��Hy-�e^�9	��L@�E�H7d8ưY�eT�w]Q�Ǘ����m)��Ԃ�T��1�о�s��_p��:�]<Z8�C�7��^���)ٸ������˘m<w��B�Y�ݽ ���e�rX�'�����p�^�Ǐ���3RQuÇ4�zyyMI�N� %|$��9O���̲Zl���5��H�l^s՜eó���n5<,x�
Վ2��U���)�h�=�(���%��s���:���ϑ�Y9���,���nm����OIi�"*9�X�Z��DM		K�uM��f1w�ܻv�����usſqq�؟1��VfY� �_�����A�	����v���k�VK��_���~��cJs*���U2 �`���"� T�/����Ad2�x'B�:\[>�����
 �e ��.v}��;�[S�U�-L�^��' �3[
�W��լ���ۊ�!>�z�������:kU�kCA�+�O��h���i���v���^-�Ȳ����i�]�v74����MKN+��5#7��R<]�.ZQp��8���j��W���I��'�b��'?�r��:{�z��m\�w�#����bUq�����>������a:���1� X>>��/s-�/�p���p �<��I�`zŮ(��c��V�n�8��k��7?��caD$��>�>|�teA +=<�&��fV�]�0�h�k�kl���)F��c�����a�ZA[���_��d���\�-Vך�j+x�<�� �����i"�c(eg��fƷ�Lc��fo�M��rwm�b���V��)�`m��@��ậ�^��j�a�'{x@+��84֣�������/$$��E>>���V\k�II�,�l��p���O��e)���Ƴ`�O�:Y��ö*4I���,�.<*xT�u�eY�q˦�F
mm�x���dR�S���N+��n�B���E{�!XK��]dW5>O>ģ�Cj�X�W�9@�ơ�4���N�ƾ@-6�#���;�4�`�:�M�}x�?�c�a�nW9�l:����*�lE�{r�UïX#5�5M��Ô���S�H�M�,�/X��Z~Lp��w\]]�>|x��[���{�s�)RDR�e'��R�V��=s�9������#����CX�n??�]�H��'k��_-a:2�2z2�lO'ڷj���3�u��u3B�|�A��0�ן�_�.���^7����ƚ�Etn>s��Y���c+���۹$	Hv�����'�?��p?�Ӭ�&�$�Upl��d��ӧ��7]�����}�� �^�tW2��(��BtM1����X"h�M#�{�9�m�}���`��[�8�w�-3ԣ|�򧓾 v��1o8D��V�#\���n'���pF̦]�1ƞ�B���Q�5��f�_��Jc� Z`�P���Ѱ�ɟ?ޖYY.ɯs��䒙*��^��1(
�n��y�S��{,���9X�Z94F���g>4f-+��d��G��FE�6�zJ+_�h��!3�^�=�E�I�ܴz�q�Rø�Vi���;������h4TTu#$�	�o,TTb �|ǹ�G �E� �|؏��!|$��y�.�[Ǯ��!\:�ɇظP.�+���d�vI�vv߅D�G>��1�Ɩ�[��IU|W��,��)�|Ê�x�{9��e��`ЕC�O�Y��_��,�c�]:Ԫlg�7*��\����⩕w�ۡ�!�x`�g���ҳ���2��eh��;.v��n?zw5�=�C��������i5@�-�����ת�Þ�_��lJ"��j+���㖼�I��~��nY���2��Ar�������lg��yOM'?����g��V��@�g���hhh�<qKKZO�w7Y�0`E�S`�Q��n/���oж0�4�VjMS��[��M1=S	~J��s*	�m=��S��N_}/��;�Ե�ںNo�$2{3�����w�����O�l�{��}�?��� �l�6� m�F���ö����������
^�$�<
�[>"���玐	�H	�z��yl���-�B�+�X�9�]�ջ� ,���mS�V�q
Q<��/!x�ش]�$�
���#������������)��TO��XZZ�Id�탏2	x6"�⑈ش�\8��[��Y �{t�bN�v�X�qY�T�(���Ĵc���4W�Ե\���-�?x���մE�}����1B��'�0_X0��G?�7��RS�SR�<���U��k��o�La>��HQ`ះj1�0F��Xn�>��{:�1�x��ݪ=h�=���8H�m��lN�a��Z�7�\ՙ����B�+M�l*W�{jv���w��N�_^0���B���ۯ��ڝՒ�������-����QЧO����B�шJ��*�ٙ?ug������jb�d�$�3	��\���Fu����Av�a�p>�JA��OvmS��M��["M%�rs�TK�ˋ�V��"Fʇ����H�-�88��Ϯ+=M��eDб�W����d�+������5�m���q����jI�����KI!����n�mkk�������Óٍh�4GY��Kϙ�O�׫7�<��_����:L�����1oi��ym&=�_�"3���Bm�V\}o�u�*��*;{p��g=c�^�x���a���誋��Z�Q���PHB�y�.K�����5� HdTTF_�E��H����z-BX��K��J���0���un�}H!� *
FDp8�_����UM��f�m���^��(V�q%s2\+ժ�(���E�DY"_����')]_����I!�b,:�����q�i�y�9m�_������p
�.�3u�f�y�?���$Ԭ%**�!�"�DUc`b"����=2�w����ªe*w����OBn�BB]�Z�������Xա�����e�����[�"�sC���PG���Ɛi�u#T�!N��B�7�N'�#3��bJ1����!�������}�_�ؖ�F��+�����8Yb�8e׸w%�b��mO�Rj�dk8��UZ֋mB��Ѯ5���<�G��.��(hh���5^�\:����r>'��$g���'��6Y�Cb�H��@�}uw�3����	_�bO��Ե �@��0S�t8�b8:�3{�;�O7kZ�yЧ�*jr�@^��MG�����X_�h>�۴E�p�se�7y���^�����h �U��[����д(+�̘>���>��v�U�j�U�fZp<�Ĥ�>��3Ev���Dw�Bz'������b�Ǫ��'i,&.�+z�����_M�o0�B�!C���W�ñ{��{�ƍ(���7a�	!a 4�#�|��+p�l��6�r&/4��f�N�z�|n��`�6L�˱�)/�?�C�b<`=I�|r�4Z���R�#���~f����r��5�\��q��n���Y� ����)�-@�2�.�fN_�~%}�F&���{�i�%�����GzU��o����3�p�5	�-�+�Nk�&���WY��J'.�5���R�)p6����+�{#I��I
�?q�޿s{5��/�"�3���0R����x-�b���UN˪&��փ�|���Y9^D�$1޸�ތ��e�}fb@�VoC*�3Vd1���E-�r�^��ja����]�ğp~�5O���P"�S�@N�l�&�y�;�\�.�5%��NN�n���4��_��)mR���I�媱���`/�d�w��ٯ��꫓&��ɔK�c�t��/`}*�_ou+V"`�\��N:���#Xi�j�j��'���f��b/`[�	TVjt�3H�_X>Q���!~�i!.��L�o|����!�/0;dblr5ew���/ ��T��m�%T��m@N�HԹ�j�Rn����;<)�RK��t`������?+��;��J�:y��9�<�Rc!<�d���f��'C&C�+��f(��U�5���r^�M��{ʹ�V՗`��&����V�l�V�[Y��M��9��	�	>ROw�(��wi;�H����U��k�ۂ]x�!gB�4n�D��pT�wE�E���G��(�k	�e�B��Z$�aKU�z��e޻!q����37��;r��*�֔�7 �%9H��T&p�{�i�	M�wF�G��ߠM��r�m�(�7qyӆt�{��EZI������O�#�C&�Ŋ!����J�j$g/�ug�=��|�`����R���4���=c�m0i3_���I����G�a�Z{?��y
<-"&��^��]��`�Ia]e�=� ��fW�3f�<)%�Z�C�V����aB���2ߟ��M+_9��Q)��fN�m�T�?A��b׻��(��~�E��WEb�l��ޕ��Ҥ��d��c
f��C�m�?�:5=]����0��ȼ�>�0�{�J6�[4v㪡�̮��W�)5u���{�D/C�T��]*+L�4c��?%�1����?��cա������joM��8����G���"��,ԙ��7�-ƜW��E��e�$�j�B���J3�щ*�d�����7ҧϓ5O p�|��t�˥��f�T�)�W��6��*��9�2���ܨ�o=	�8!|9E�Ϣ�r��gh*�+����N˷��p
Uwʢ� �դ}Qα�O/��D�(����{�!�v�W1��'n���  �9oN�q[8������hb!u��j{��\DJ�_۸{T)f����2_4�{�1V.���ֽ;���xd�%�ݰ�C���Ar��O�ה�!w�=������}YGl
�K�r�f����m���\Ok�`�h��x������vN]]��C%��@2;�ٿ{mB>��0-c�˚@ ����|�>��E�ׅ��`HJ�M���W��x^Й��T����8n0'u.RJ������( ~ �~C��Һ-��h:�u`�8	���o!�x�eJ��-�R-��eCUZ��eR�J��͓��0%b�z���X���$�m؟�,@��D����k��Z9׹�B���XLt�#�k�Vc�V�S�[���CbGY
�k�6J�?W��z4u�T6�(�H�C��o��=88��{�}vc�ɣ��Ú�?�=���BGy��[럅:�	*;*+��ZV_V�|\��p+�	�q��X����ic�՘�gn 4�P
��:��L����G���@�1�ɖ���E��(�S>�U���m�~�nRA��e�__Y�x����d�k@�.���������U���ߎs,��eb���]�gbޖ��>r}�:�8=a;��{��p�2�L�n��q�@�e������=����g������� *�<��uD�U{��Cɛ-IR�BD4u<��-�������5�Ĵ�N��ij]Z$�B)�fq�5]6f[��O��~Ӄ��	#�Pmml���U֒8�a1�l�U��K��*��@��MLL*i��׶���F��`I8��[g�[w��KV��#��2q���\�n[Z|��E�_y��s��w�+���#��֧�#���W�6�Ҡ�tO�iXʪ��b}���x*�e�J�tŽ[��ne���b���8��������LGfO��r�ͬ�I�eG�:��nK��&-��-F���I#�(�TÅ��Ѹ�@��.=e��Q�Pʧ�,{1�g�-;w�1�������k)�E�[�w�=7S5�-ev�г���;�P���@�r�Sq8͸�@���O���e!�LxԪLi��
�[���HC���_�����9��!�odh �[�ꟽ�9	��uݭ<>�k���Ac�`�ϗ}'��=�ۮ?��9�v�kd�"\:��q��A +h.]�5�t���b��Yҩ�fN��&㙌e�l˲T���[��N��R?	�'�=����2����G�K�q��[����-���BF�6�,�\��
3u�4Igٌ���ie��&-�Va�ϼ�j�]�onm��Z�!j�8�N�&k��ܜ��Ⱦ�e��{�p�&�p�����)H�a!�Dk,n�����igKJ�l��(�f��*��v:�V�5���8�Ԥd�pm]��NG�f7��{��5K�� P�����D����a�����T��.L�i�cVi��$���,x/,x����߄��D�BIvLF�(17�"�,����͉����ɍ;ԟHt8I�PQ5
�*�$�q�"�6�/ϥ�Z@�n��ͨ�u��fXJ�L�S�I�ů��zΝ�9^�A`���F�ش��F�$�ה�����~`����JV�&D�2p�w)TM�m�f�r��X�|��I+\J5	�����7�box�\��ޠ"����]Н0V� ���Zrgh^�UJ�����P�c�*{�$�"�⤿�*�9e�6��bY�`��j �|o/$�����[!��8U�&T-�8ֈB�x|H-�rtF�UL�C��VKJj�Ɂ7}�Y�^��z��q߂�Cz�u�RBʩ��馋�H]lN��]�y�=h��x��������;�?�PX�R��Rv˰B��$�d{
��X�f�	`T�_]UL����d����ts19b�/�e*:ک�`�d1�^?�:�t�m���!������ң����v�+�����v��VF���5~Y`A�A�#޹h��W�VE�ٛ<�����BQ��>�h���>�����r��X�l��~"����;A��Ҫ��
h̬��k�m���k�)����fK��G��Ī�N�̡�]�Ն'�n)�C��Y:}��m�s���#�$)�����s����y����u�¢ ��aH-��ٌ��n�L�O���l�� ��|������*hb�dgq��o��a�]�q���v� �P���Y�s�6~���'t�6�ki�?��:����U$��P��n$������
J
H���t�Ơ;�C��c÷�G�s���>�~����s�5���c�9���7��ݍ�a鷼�3fbF9r%��7ͥ��Z�Bq�+R(�	��+uYV�ţ��]��L����Ⱦ��oΔt�'/,%���E�)v�ojn�H��U�1�C�pC�&�F��R�l���$4�L{7�6ħ����b��.��ȋ�PsW��v!0e�_#��]�Έ��0�J����<�Q4����A�$)U���j�#f����w��R�畴}��ktE��bl.�b�y=���gʏ����Հ>�ȿL�?*��&��s��iW46�1<��5�˲�֟��f������m]k1)�n�)_0]H�\����̎Wrٔ���Ï�� L��ا"�7㽵1���'��g5�1b���g�P!d�����j�#��b4eAt�¥��-7��KC���@(g��Q�p��3~��ɞ��� �_1T@R,��tv�a�k��e);��u�=�f��X�$M"���8�{Nv�� 2�ʨ��
??�Z b��V�^u\l�{����Z���{x	3.����䕃�jꏔ�/����{�^g���\��ͫQ2�C[�p�)�&w��iO�ЂY�{.���I�?���]ە��q={`ji�6�J�{R���d��T��������U�qL戨ӱ�tTǗE6Ġ/������ώ4��-vC�6M7z���̣���Ѕ��o�K=-�h9X�iE�s1z��E]�����a�ۼD{�W�Q%iz���# dӼ3���Gܹ�9�&]����	y;Vw����M���y� �(�f�tGg�t�WS~��Z� +O�F'.�IS�%�]�X	*�|}�%��U�UXD��Dv]o��}�zn�"�N�7�K|$�7{Zo�fњ����jEk����	���.�N�����Y�rם{{GH;�b�N��0ƕ��N�~۱�s�]��"A5��O#(�1&����+����\Xy/dH||����Ϋ�T�į���'��u�eo��.�7���|nT�w����ff�^����C�v�2\}5�I��WZz����(]Hl�!;��E�b�>5���f���a����9�;v�G+O��;t�ʽ���/pD qZ�`2v��{�r��}hĠ��+�x����5�����fqeś̞�l�/����J���18L�U;�7B�4�\� ��n�,����ﮒ""�}W\�3,Ŏ.�Z��w#����-��ٹ�6:aL�2  u^�}����2@�WBy�CïHsR�q��n�B��P��v�������`~�Ar��0�Dk�:o��[�s�����z�./�����3����������q���w�uįL۔W=r�[��N�pZ�.�-AǍ�@.U�P���=��H�M=H����2�ˎ#㣕ykrD%_�[�\B��vw�܌�l=�V���^Nq�fL�3��i�<�C��::.��&j��N9礵����i��O�̷7'Z��<�-v��H��l���R��=y�!�㫎C)wLu��
�g_~h��ƠA��#B��2��K���"�:����*=�P�v#�
����.��"y.�@� �~ވ|�z�,Q���ʚp�u�j�`Uj�<���<��ޙQT<��B��yF����j���ER9`�	�f�ۍ�7�
��V�Ze.�k�E9�w�[*>N2�**e�x3/S�.Q~��UY��M���KKgx�"���K"�z}6r�*��+5�zZT��R|%�nTr��Y�T�?@�(�_W�2�44''cJp]Zi0)j?�P��@�e3;�>��o뺎��;y *My��3�Dd�	Y�����An����{.� ss]�\�^�z.�����F�A|g���iwe�־���H�W�2��=�:�]��hm��&z[�`9�b�����Ⱋ���\L,z��J����EO�@�(�Ӣ��&��qo疅dkf�@�%X�ډ�j��I�oNHI=��i����m��ͪ�E�v���c7�8��z���ǻu���'���-�x�pv�n�qaIX�]Z�1o"����_e������IJS.�{^p��3=��7�֋%�]�֏��R$2�_EJ���"��+�llt��!b�j���fZ�&����uN�h���zXu����5B��#�'55{�C���[�s�����~'�І&�����G�\����A�})�=��"c=����K�
��.���C��$^�m�O�N~ؘF��X_�h��sc��g��Iã8vWڢ��%|�sۣ�~���o�E�����.���[�jt�d|1�yN�_z�|��w➊�R��r�;�0��׾+~���9�lli�ú�h7V�w5C��3��/<>�^�m��K <�U4����zR�*[���K�q��2�r�)��^Y�q���2�o��B{��y#=ڒ��=M��-���K�I�t���^����?'=�fـirR��-���� �����',--��ΞPJ�dxa�,�����)v�ZD\��B�V��L����Q"C�"L���z߿ƙ5y�M��ut-6�3�hK쟻��bj��e�^��:��ť��kW�Lg  ��i��%\쯜�%K��J�<��<v�ªx�S2��#�7y�_?'���?<::z�c�6T��А#��[2\ZL˱:�˘� �sV�����uٮ���f��t�\踰�5�ڰъ��]��e]6WZ�K��)q�p�O~�y�a�VI;[G���W\A�[s���~���Ą:B5��{bFƆ���{�m�)�����_����.nLz:�5� �j]K�hl\��ZE,o<�g�x($N�������Q��Mme�7����ߥ����M�rbh�5p66O����t,S���
��R>�����F]�C#�"��a(�����K��׵�F����zU�e- y~f��1��P���D��{���H�իW�4�C�Q�o�ُ����C����~w)��yX*ƿ���4aNB M������Z�E�޳j(%#��N�2+����Do��-l�wD��p����>g+d+�YLL��(������'ś]*?�9�G��ހ�M���9^���GP�g���֦ވKJ��A�VW'Y�UE�$B�T"�\~2؁��Ml��G�oZ�?��}�ڎ�R9gf�Ar���V��N7&��}��Uq J�G��j�EF�n�9�owǵRS��%����<�k�����Zf����E�o/$ؑI�ʽ�p �4�J�T!����8�M{ c�ڻ<q���hL;�����i�d���h��Fw��7/[W�|��n.�!��W*�E�E�?���i�5X���.y��7U���h-đ��)��\�wt�Եj�n�0�^�&���R��c/�`MƜ�)i�B9yy����f/Vԕ�'1a.�y���YG"e�x�@� �o�Xe� =�}��u��g�:~���b;Q�Xd9��%��]��2�8�����	�R������pK�e�Td���£li�Vޣ������GT7E��Y�qvv��v��`!0�=��݁.QhOqKk/-i�V�+6�`=���.���Ɓ��^�3p���vc��-M�ӎ�����&ۂ�����͇3�H|�����Ǐ�1�;w��f�d؈m�Dԏ� 1w��_߁�������ˑ�Y����5��=Xx��W������!�[�T�l�o��zw��I�Dϒ����3���|���d0Ŗ�8�?�LS��jb�ZS���@[�ڭ���K�z��Ja� ja(*��)��3�
�ɲoN�wNR�m��b�bCX�g���$f)����զ��~b�����E�a \����0�G%�<P2�(G��]�J"=� �?�h�����b�*�ij��͖^B@H�Yʁb�F���g�^��P���f���h5���Py"c�����t�%F]���5�9)�&��Ldy,/-usE�u �?�j:`�1ш񍯉�a��o�*�mv�G�,n�ul[��(m���/ˍk�N���W�خlv��nz�O��I��i�f!��{n�ro �	}�]�
b�5I%����.�\ވ�M}7->�!���h`�m�k���te��m�dP�������lP�c��� �
�=	t���[���R���T;���M�@� ��A�t����/ڳ����z��b23o޿_N���� ��UA�������6DY��:����F4Î���n%�mX�K�iiA��>$�|~�kU|�h���V0M?�J��Q���i3�dI۾}�kY�Z���{-�B��Ϭ+v�A7�`d�A~��:Ղ�0����׆�@`�x�G�S���Y���I�SR��|�������J�s�'�}�|����@M!�GDh�L�XQQ���|3����T�tn�L���7zdat7-�J��$P��^b&ݻW3�%��.�$����ܘ�{P���|��͕���^ە�VND���%� ��3�_�ϟ�V�`}%h���񶲲2 �;���S�K\h���О�<&��i)��^&ώ��iY��P6[k:��y��|3C�����N���C��놶���Ö�-O#��y\7LSF�t����*��w�C��'s���k���ӝ6��}V\�Y,�zzD	d�La�f�_���t�DG�W�����`�����D�)�4�s�H5S�isX�O�x�V!ͩ�x����,�����jgqKs���� o�@/5�mS�]\0���Q{=�����t-R��\�ж���@�0 !���W�� ���6�	9�7&8�m:zt�	����?XHer�o�0����Ė�����CQ�s/x]���,��k��W�nx+K�V�u�Q���/�	/.(_X��8,D�	`�s�<�.R�x*�X���˨=�(�� F�?"'!�����Y�������W���/��4_��K@��}M�R��-�M$��ea:�ڵ�NAK��]0lh�u�p��zA�ѹaecR���>�Z����yu��Ą��݇ �M㈳�z����NZH&���'ERr����#RR*�3�q�ۣL�1t�#��&.�j蟟�0����h&>'��5���4f���β9B5�������y��XAAc��z$��Mf��#Rtr2u>"Ĭ!k����G�ך�.Q�=otc�RS�7Tf�%��t��>�0e~vq6�#�_��n��YZ�^�
y�)�E|m3��ePY}f7Q�Y�#�v�H��mng+2c�C�����~چh�޵c-��m�4�G�`L���%��3��������EH��9[ UZV��8[�(�7cЃ��Lw{ ۗZH�[a�)���!az�ڨ|Z���XPB%۴qkܜ�y�˶����
߁�M�uq�m�X�`���=G�-7"�����_g���ST��>(f�fR��xXڻ%SP�����Ԅ����J���z{D����jEذ��Q��ٳZw�� �!#'�hpM����bLF�3߳^��� ��hٴ�/�y6=�
��T�߫Jx���s�x����&{&4�(�\�J�k�����S6WSS۱��T�5H�H�&�[o&(���ʾ@3�C�S���hn"n�YL8��C�X�--�))��eO����T/�"��k2�P�yuT�pX|ڄ�R� ��x���6�g�gy^�B���;���M[�3�V⪗��.��$0DЕk'WV��^t4͵U.\�S~�������@.�9#�3L1�S���g����?Cǻh)[v"
����,�0�vEʻ�8ׯ_w���h�P�Nîf�@�˄�z��WB���q^��('S�9ݶfp���edhc�h�7<�U��굼�4�=�/p��h]�k]��]��74�^"B>,'�������-�8����&'{�����ˈ=�Yt�X�$%%�+,䢦��NZ����b�eg�GD,�	j�< C�P�"x����<��n���Q��|~n���)�D�1��� ЭR
V��!�r��..�����9�q�1�a���c��h� �B�w�rs�V]�sF���l�-|R�_���b�� N=�u˧���U���Y��')�#�@������v�#3Ļ�^���[��0�-vT�K`z��vC��7�b�Q|9�]
�$���{Ϲ�Y��e*5f�R�®�v�-�g$A�  $�d�q��eP{s�C�F����w�����TTT�"/� �u*�9c5�����7ݓ[O+����n�k@9Ș)f��i7���I�r���<�e�F�[����]߻	V�8�mWn�8�z&���w����Ƕ_�{\e��C&�1h�HE��B��@�|�FXHH$G����5�gϞI������m� �и;w��W�g��E���6����Q��2�iK�����0���y��u�pw͏��\��;M����G.j.D���n�rAe"���9�ڞ�J�������"���C��� �fae�#$���1�۶G�??C���a�M0F(` Q�Y�� 0��+�Kjkka��΢zU�T��q��|���gX۝/�ۯ{�����0�3O��FUlW�]S�et�Jg�^����"�yaʁ�}:��C�=.d`�gg��a��MpQ��zUʼqz�����Cf�\�8������3�!�S[[���o@8���fz�����������
g���*�Zl~�ݓ���Oo"�`�XԱV~���P���].Z�Km�����)#�v��u���/��m�y�K�9b~;�;��N3�Q���q�zQ����A7Z��]���Gd�+���$��~���g��9��Y)� ����|^3�CD�L�,��#R����Ҕ+��o$�A,\�g��%�����X:�N�Oe��"-�P�Y�H��=*���
�^��;��%�ƙ�wa�Oqf���!U
ͫl����{�p�� /��Kwş�_��K]�'��zt1�&|t�MD���ךz{��t뽺���D)g�TG>�xUv
瞛55�C@��<�AH<]h�CP� ��K�9�����s�C�r��	弍���z�:����D$/�=XYj��>\1n:�Y_�!����f2*��ĉn'����_A(//xZJ����<�!rOLP�S;c:��0>������q���	�u  ��H�?J�7�'f���)�8$,.M]��a�C���X��ִv�GE� ~�%@B��A�f�a�n���d�ғރ��	����յ�s��F;e)��k���wL+�r��Ś+�3����k��M������������/����������L#UT��j�Ol�3�Ą	�,﯆ }9��S�c^A���$zG{g�It�2	���}W�M��6���"�_���V�+�<����c�fp�>��h�Z�j��W�^ݶ�^��Q�|����LB;��~
\�~B��rk��З՞7�on���B���o6)�����]��x���?��?�0-�5�z�Gt�)�P���?L>�]�M��J���s��hF W:�P^!��v̢I*4�Ip��z�4O��[+b�C<�ν>'w`��7��zm��23kg���hظ��n�+�>�Hr�MD�r�
"�Jꓽ��Դ����A�;Xh����E}�z�)��-�a�:X����b�C��R+C�٤|�1��+������"]���P�����N^���=1)�3L_�u��Eb���B�%=?o��\ �U�4�|<d�貰�����S��^JE���k�[	�t�m����*\�§�q���%�����;��_������$8884_@�^�L����x��@��p2U��Rͼ�=x]�E���r�G;'�J�h���3�$����R�Ǳ�81�`.W|f/�MC;,�@ |׳u/��@���3��3(@"c�q׸�O|��,�-)��:�i��?♹�9�H�����Z;�\F6:���<�&���=���\,{ɡ���yH� �A@X8�`!p�ڎMvN^JX��!m�EYo�%J��1�<"���l�Ml
{^��t�.>4�*I@;<4jJ�S��!�����z&s��uO�����W��}E@BB�RS+�y*`v�\hn�9-a��]к�L�h�8�~=��C��鸐��v}SSu��ěxD�UU�T�F�L��2�o�(Y�NAN��,�j׎�Ru�PQ_L�Ee���P�2"���ޜ�<�\꣯q���������z f�����������U�2�9ѻ�����64bЀ1�M]�̷��\�cDH��6� �(X�;�ތ�Ok�F���B�  �RSşA?�>�}�j���� �jxx���j��
hjj�
����M4�j}~1�i9���M+�6��ISH��5j|R�j�_��i�������mNN���u�а��o��z�:�7���}�8ozy{� �^C ��r��4����$­�&z�|�di+C�۬ࡍ��2���> !Ԙ���?Z=�G��1=s���N>8H�)?��*{ߤL̇T8[eeq�] ۊ��ǖT�,��n��A#�4�^� Fd���z��� *���:/Ұ�%.�yu���߇�K:>���������vjze�M�K�/��#��H���|����J����
��@�MGh��� 檋WZD9���hi}233e6jAS�
 hM]��.CR�l� �k����������>W��(ݵ /��I�RH�J���ꃅc$���Hx����%@���ɟ/�~�sNf�CZS[�}gCTGGg�z��l)�^~_��8�m���{��i 
`�f����_��d�!ಚ Bs��Ȫ��QSS���H��1��HM����!���j��9a�j��� 	xZ�Ă��ʻ�ӃK?fxի�D/^o�І���q��M%��m.��;��w�����F5�q@ݮ���o�XPl�s���NZY�旡��$|���ɣ�
�&��D~��UUKnb `���[%���ɶ]�9P�����=��9��Z�'��?ۻ/����&�<d�@u�����!���dUHoIc>�2t{�Ɏ^�-Hzy6)��[��ͫ�e��d>|�z~F��94r��hdh��f39�%E�͗�c5f�r���,G��ku��a�_��]	�_�/��aֆ��a:e0D�mzzZ����x����o���h*��`�C�*�#4X1��y�g�M�?���( .)|;��?F�!�M��2��orb���b�]8��/�/hQR����F3 �/te	��b�A
n{O4���ܠ޾FJE.k�
^ss
"�������.#���/���rqR'Jy��'Jy��'J��R��"ػ�rߍ����E;���{���1::��{�V��4�<��7����l�'���K����Τ�����@A��_��~�����u�)��4#I�� '�������(�B��[�� ��		A��w�z~lN��p�J�>W7K'5Ä|B����F2RQ�{�*�>��;!���	l��ǣT�ΰ[�6w��Ep�3` ��g�:N�F�$o����@*�1 t �ק	h�C����32˝M{�=�'E��#咭u�V)�_����:R4�����x8�uӺ�)G���D�ɬ�dt�]=|��y�}d��n,��R(���g�Q<aY>o�e;Kg; 7&��~����̌�.77��~i�v�xt�ӊ����	ab�]^�EmL���S�{�@LBl3���v���P	�͑�������۷>QH�ަR�K§�ЌLM����y�^��#�ߥ\6)�w�:��w��#���V��Q��a��;��a�ξ�s��ʤ�����ֽfvu����g�)����C5�bMN5�͖z܏}.�A������)nUb�+g� 1P���?�i�\�5 �ň����wr�<�Rbw��o-����i�5��)@'���H�E2&�%�����R 	����A�V����Ӡ�/.Q��O#��)unw��H_�(*(*���]�j�]��竃�F��!v�� �����-W���B�EU���x�i}XB�0�5�g�B�̗�,�(	�{�/�7خ��24$I	2eZ�_�b�<}�Vc2.���l)�^wTh���F�1�{}>��"63���q-7,H ��5��/���"7ZYd6�9�R"ʩ�� �]V�د�-c���u���-�'�E�F�嬲������떢ج�q�߿�5���<�����Q�w�-I��w�]�bԃ�q�{����1��y�O�P��!<:r�x}���PXVيPkl�~�l�!��k�ڮ�!-�@�33�lkkk�筸��\�]m2 8�l6f��k�?6�֩k҈�Q��}��5�c��hj7�M׳�a3�j�ΕWlG �R�l1=?3Sl��>T�T��C�C�)��<\d.�V��uֆ;[)+�F䗌"��W����)j`a3��.4����÷9aJ�[!L5�!��\���g�^^�t�_#	�/qju���G��%4Nj/u������I8OI7�:�}���-}�ݵ��PF���沦��1���(?�$&�`����B��J���a��� Cؔ<t�@�C���t�b	>����[
�(�$q�6��cs�H5�[��̰'��()�M@o��f��{���"C����~X�}eL�8���#...==�l�r�rt��؎������X�bȳ��擆mg~�z���9��f��dgǥn�ԥ�:�����;�����g��ش�E����K_����d]�[�j|z�=_79�����7����V�9���M���BV~�5!�9-u�m�uq�Y�6��F�]C������u��o���	��O+��r��kzz�ؔ���<5>�Z�4���h���`����ǖ��s�s����+S�.~ə��tk@z����7:��;�W}I�(�Y�<]�
u\����/�9�p�GUn`xqc,�yְ��7<l�W�-��;���
൴tT�g3rr���0��py�� �ќ6���E�dK�I/*H�)n��#cz
���$�����J�ĳ~	G�J
BBk��d���=F��q��^S���q(.6sb�
��w�Bp7�=F3i��y归��D��(�;KVVb�Po���	D
��:��Z>춲o�bA�T�$����=�l�	��r�#E9@��n��/�H�(�i�3d!�5�y�l/t�9On��z�1��1P����ln绰��9�e��9�=�� Q��w�a�����ѵp�	A�Ўӧ��h����ÿґRQ��&��4D M���]�#��=�	�_?p[�1X���Ae���}�����^7����98��O��Hp����頾j����~ ��0x���㬻�a�M庼y9rN�8��`2y�x���Ծ�lޟ�c!��w33�k�<8,�Q�-mS~aN�e�s8�3n����-=�8p����~	9Vpc���+�Ó��W��E��O��?��H�AV��a��$jv%�T���
�$zy��������hG��u��9�`�&1ɂ��ϸv���*ބ��±'#�R>G1��^^�q'�7k2��}���>7�'�d��@2�P`y����UgGh$Q,LL
1�sP�ʤ�e��267QV1N�m_��3,U4����8 ��\^6����lR]�^]�'�Oq��?k��n�2�`{�:�FY���|�?��0�����'�u�����X�tp�2�1��)���8���x��t�Vq|v�;W��s�`�Z8�ؗ��V��%)h�:&k�n'������̶�%<m1��
s��CR���q������[Z�%��G����5X�/z�?�J��ӁQ��H�)0�;ݕ�E>�u�?��F�|~�}�萖"yV�=�ؓG�<~����R:�Zf{���|b�Zb�zkى����Q�
�Y$��6�r�}s7�fE2�� �����g� B@��{�컦����^-����u�Z��M���n�����p��o�ٰ���k4l�zO��˾EF�� ��ۛ�lb\���ܾ��/}��\cH"|��S�{<���S���Z`J�6�:���t��`�JFJ5F���U�0v-n��Z9ʅbcb[����/�|���s�p��z�ʑ�T����3v�gC�E�m��v��*���#���[���1R�?E�T���2l��1�X��Q]�W��2��{��@���~k�W�-���Q����.�{HrQ
h��j>َ�G���W ~�7,�v?�_G�R�{:�݇EMstű ��j:�k�#3��]��g�|�	{�\�!@C�Jl��o����Yݷ���#E���:�Dx�%HN��MI������TA�R��>�>�[*��ݟF�>������i!EH�O�xMK4"�~dˊ��q����g�������,���aw,�eq��ݦ�+�]�0e��>:� D��H�{_}��n����.RQM�#���:0�m�Ⱦ'a�eTO����Lr>j0?dd��T�� &\���J��z�[u���s��{��oN�S�X���L唗=z���VҰ+������59����j�	Y�� TPI��oT���R r6�i��{�31�lH� Sk��n�1�_�8�a�k���JG�ΔP��1��w>ab>���ћG�=b.@�v�ﻏ��򘓖7K���#>)2�91�߇ i���y]~qd�)Gି��A��Ǔ����=3�AMJUѸ�(1�C��TϾ�΃)j�.x5@��y"��N	_�>_���N���®�Țz��B�� {�iߚ��c �=���	{���  ]�:��s��Qqg�UҼ�c��b��~�/Ggid����5�=��L�ߗ*��]e�*�f*�Ы|�#/�<W)�̾���O�q?y����%ryre��t����ߧQ�&
vdCh��GěS�Ǩ ϩ ��wn�c��Ϸ��l,/??��� ��R�w9��%�="��1]~���;#{蛀�s�A��/�����M���ޑ�^'$ Y���۾/PӮ���v�����v��k�,�ß�-|kY���ǡ�4�,�~DZ�n��!q$t�FI�;�n���)�@�Ѯ�}��>���r�og=��N���� �w�w$�������5P�l5W�U���g���<E-7���7lu��K��X�;"<��=�$%����M�$?��{���(K��#��2
@������e5�4��]q�,P����3�q��$�Z�s��M�;�G�%kzS���GT#1;��;٠�.#����99�ǁy�;:=˭��̻(���Gw��̀P�����m�G�ZC&o������e���d5Ӈ�|��{i���Yau��L*K(L=S��ϸ�!9(���h����L�4�O%ݧ����ɚ���9":X�<��x�w��k�Xv����ކH�ca2H6܃�<�Sc��$do�R&z��\"?��$��u><ت2MG����fo� ����ʃ鐿(�3R�x���'��	�徣B$�`ƪҳJ�ޯ�?������iD�=�D�j��^��0��{6m�1�4��)U�Hӡ �|{�9�@�	�<B.��7}MG��C8�y��m�}�����H�L�Q&�ݑ��I����O����:�����9;��X�d��5����ine��	_�̊ΦL�Y@����ۯE�����[p������T!+vc�9v(GňL'���_(l��]�"B�K�G���i�*)���=~6B˴�#��'V��w��)d�K__�����#iRj��I��f�6�Z	�Q�=�|�c`r��&������L�$�c��A�\+p�T�o���({2��b��zT�^�	��ŧF�1~E�.Ft�t��ά�ꑧ�H����y��}E���}W���o�?��L���F9����i���hup��p9��a��k#��=WQ�ߟ�y�\*��(z�Ȓ��%\)T��Ix�9�lX�Qv��@JU���G�n������u���q�Uu�6)��`�C�P���j�Q�s�ކGw�R������?��x�^<-�G�Q������"c<�\��)ǧ�u� &�u�����	,�0�O�f��}�F�5n����� !a��Y��N4.9���d�WA*���1�j�����#���1�,�{j��/�#��{���⺌G�&rJR*��`B8�
���\&�E��Ȉ����4�.ab_�X��yW?����@�������a+���4B5����(2+�� H�0��mn�oQJ��{��i�����%�~<�ۈ�rjƆ
Mصi��G~;����^��#��E��E��zO�O�|���~6�#V�ĥ
�C�r�_WA����G�r L�)xG���z�q���1	��8��&`\tbGOvh���$2��U�h.�,�럓\'J�o�]��m��e��S�]����h��D}�
o>��H#�K�� �Մd���������/�� ����Dg�Ñ����҉�0Ľ3(����RMYؙ�Oqq�����{�o�I�bQ����6Ot�cs�O����Xi����_��x��'f8Z�&"v�Hmo���$�%Z�a8� Oy"�A��D�'�<� Oy"�A��D�'�<� Oy"�A��D�'��� V;��p"��<�����лQ��1j���~a�.�����N��7�2E '�@����}�ؒCJ\�vo�gF�ē����������v��_ԏA��D�'�<� Oy"�A��D�'�<� Oy"�A��T�|5l�ie)�y5wK<�yf��`�]��}�N�Z��5|>AF��2�Ŀ����X����l��7[�oq�o�5���5e��hs�4�JDT1A�:염pJ_�h�Ry���X�Qb��=yv����NqQ��E�#<�NA�MZ`�3t5�J�w��|j�E�Ҋ2'��c�nk�F�l����[{���8b�����L�0�]񲝢�w�p��\c���P<�|����Z�6���C���9��Q����X�at��^��o��J��wa4:ή�+�=�s_F<MS��0�/M�P�԰ix*�����pTJF��sYV��v�.}㺖��f3����a&�� �{	��{�k�%�����!p����k���1�9���Ll3��> ��D�ag��#��|��H�hm�38�m`ȸ�9���%�uF~������8�d�S���;�{?y��i�<[!��V��`����}�"�Z3�'/�.��۷��ܵ��;���*�����������.ő��� -({�㴺"_�8��С�������!(�9��='3K�L�U(�R���:���[`[Aܚ
���,�9�W!����}-�_g����PQ�=�86�i�!j0�5��2E��u�S�;�@И�B���J�8o���ƥ���l��v���Q��Y^l�����<0n�0������r�f�����CG����Uz��b��u�f'10�|Pv�d�>���Yd��Bȝ	~�?�)�� ��d����T7p�Wd�|tk���x}7 s �x:���� t遬MG5�B?r'�]7�D@	���_��׽���GK>�G]'�����	�����S�d���e��z������\�����p�t(t~�8�	.��_aZ�YnS��������1�N�Un{^M�*�5G������/xi�z"""F"���ngE��e���R�+�>��k�Ou�[�QE��ͯ�\�P�$'�8>)F79U��+Q�ק���PJa���`܆��{��y�S.�����˛艹��{��_2U��aJM���p	B���~/Ȣȱ���E�짵ki�G���I�k&�Q�x:�Db��i���k����H!͛.��̩���(��}�}҄�~��a7 IG��4;���f�[�4��]����D���,���D��<��l�2�t���T���e�=���!�O|���.,��
�����PJaٖ=k��:�`S���~W��P��l��9?ٯ�;�����:�a���u��h*� ����j��;�pўUt���G�cq�����:hR���;T�Rg���c��Fj(k�]���/����.����wX��%�BV��y��>i,�ĦrV4�ʍ�*�fu\	G�O�=�֙����2iu���eAo�L��	��E�?�܏ta�b������q�<�L�����حw���^��z��8�J�+����vԻ���������m.�RS��{�j��+6���������0-uџi�,FZ��=����.�<����h?ki_<y˽�a/`<�罵��䧳�Y���8�t�9&��T�01I���lSt��b�/�J����*)Q�p�[r�Nɣ�q&ؓQ-�z5��� �ƦV��)�]'�>����{%EE�!!!sWV{cU�ƨ��2�&3�\ry������&C�f/Yu�V�sfuk:�U��uo~�uƟ�¿%�W��]gc�=M�t���:v>�aX���ZpFC��T���g��qݎc��0 ��oL�z��+�Ͳ6������#���~ؗ���=M���*�םͭ�����n����ym\\v�Ԝ˿�/Y^��]Nd2|�K8Q9E�d�_�^���|W���lN�̀�|�3
�/Nf	�	�(+PYq�	�㾛����]�cO��?|)C�yC�S,�g�-�\7LPvh=�Z�-U�Isٸ�$�}�mU�k����SU��wb�Lltj��ysw[D`�}�,�Ӆy��o�w'�o��;O75:w�U �4�z�~ݥ�A1f�-s�iOr�悟4�%Q�A�:mZ��c�q����M#w����h��j��O���Sݶ���r�#���yǜ�`���yGtt28�ħ�$��F�F�n�N��D�|�
���w!�D�4�a�!�C��vm���{���}=|��W�����豧P80:}����Ǻ²�]my%�����P���;Lx��x�N�N�ߨ���}a�1�<����g�F_�E��RR�z��T�4V�w�w�"^7�����sGd����c�Ǐ�|�s5�/.>����,�Eŷo�HT�.��JV��wa�R(�]]]�)�w6�^3�n�G32D��n�llmk?�5iť�6��6Hr�����#!����|��e��RF}_nЕ^*HAA��dK��gt�27=~���:�I���� ����zE�%��DFמc�}��"詄�)pmT�@$\��ܡ;*,����ōz�3��n������s����@����S}ձ���O��^?i�A��|��R�ؒ�sTw�
cq�����c����p/��	�����⇎i&&����ʭ��V�Z4wt�W畮��)����U洋�WM���Kfݺ�^\�N�O�����+��iAMͷ�=F�������� ;D��)��Y�ɩ)���9*�����b?O�3���|O�.����i��������~X{�bh���1L�f���^M�`�5ˑ�M|""roR�!���n�*=�����>�I��FJי#�6\��dM=i*��ŵ�b�L��7 l��ȘY����8:u���g�c-�������K�B�=<<��P�~];f�Y�ġ�8'|e�v�ϟ���ڮ�HH4�a\���\4_�,m�X�]�o@��ć�����!�9��%q\���!&��t���n��d�~�P]��Lr�OV�ξ�U�rww����ab��w�U���ySW��2���t�˰Ż�i{�*��A�x�YA[,�|���>}���^N�F��n/�%{y��]3�{t�vO�s����	t�������B�[�u~$�*p� .*$$$E����^C@���ԩ���ȼ��Z"�!W�����P�W���8���pnjj�6��i�o�1 �˶��cc���Ocyq�~¹���[˃��l�L�b�(xf�T���y���2�vR*�-�N������5000�j%5�O���w��htP�oV;�)}J�NX���B���@_a=2�p�	O��q\�D�r�2~ɰw��J��B<��{	�~9+��MM����5�����dM9�3]ܑ���D�n�98:fUzbA�q}��h�k����M��v7"��-33Fddd��ʂ\q%��G�� بY���F����ͭ�AHU����8�(�����9����py%�(s@�3���9[O��RL��z/|O�O�W���!����=��i�*�r�m�Y�4�ǩ�>3o}�~'Q�qz�"�5���Nig��zߦ�NL��v�fg=�?��e@T��6|���
J
*�)�5��tw
"%��ȍH+H�R��1�tw�  ]C� 󜃿������_p�4�9g��ֵ�k��I���?���+�}!J!Q꺙��߳R���u���?BX3�+�+���ɡ�����ň��].~~�W�~��U��<�����`�w�刡$���+F��ޞח~_��G��&�7������q�kтj�&$.i��o�+w�������l�B�/w�=�߼��� Y��b�k.Dc$�����뿑P��J�>9
`0`$��^��,�㵯���b�}	ѧ���@ǀ&��I�O����~��Ni�n��#{�����/��)�{�����{Jп�9�Cfc�222�!u���lGhj��QH��5�v���ؒ�[/��)p��+�]����/�>nWwwsW�1�b-�:H?p���t��AGH�� \��W��I��3GGǄ-�t.<�~?Ҵ7-m�nq�v�^M�&������Ú�xw�Q�S�ѦI��`!�*n�m�7����Ȑ@\x����ŋm�jM�����RH0'�Q��͏�;Ia������U��1A(�H=�arnD�M�r��I��;Q��Ц��4"?~��8����0m1rC�>��HF(�a�DO�	Z��4���1�a�K��xdX�k�W�M�L�~�U��Hm�Ј�i 2����zlz(�'uΛ�f����Ht���.��� �
��ee����#�bB���^�w�D�y��Fھk{S������ґ��8��,JcS?u<J�W�,m��� "�L�׭v�#e�l��c5.�@6�	�r��J�0`��_Y��Y�q���x�
�n�P.��f�kY����C�r��b���h���@�����}&&&�I�٤2{�fٷ��v;�CߴX�n~���H��#��*=�t���Q��x�������;�������R%�)�:�\��oݏh4Q����2F�.E�+_�q|+�Wτmg��6�g�;��=��UȻ�LZ������@iGE<BԻ��EZ�5AM>}�@��Y�X�c%�W���]0��@q�o�C�{50�n�E�Q�
�\��L���Gl��_���B������@�H��>Ƽ.�n.��:�I���Jɘ�+�$-��I،	bƤ�QR�MCr1zW`�[r�����|�xn��Z	�(9Oz]���RCcU����06}6����CՔ����x��`�� �����Ѫ	p๥�����������}iw-A������8�K&:�R�2>>_zM�d�jj���l�p�(��qek+�굛O�"W67��/�@|�LJt<A=Dȿ)��#K�LڣG��s�U>��H?�jg����o�e�y��c�� ����G�O������V���b�
�a�f���ͻ�4A�u�ӎ����~�+>d�ԯP�Ϊ'/w�=�
c��F<y	���X�(��%�����2����/�I4��ܻ�����U��.�a��K�n�J���7�d���f;h��K�c �ѓ�]�4o(	�e�#a��\u ��F4�T��v�{g��}� ��^�BL^���l����7Pӕ��D<��b��K���c>;;��Tj ���H`�kEt�ڔgX�ï?w�ʽN@�1iZ�����&�0y�_[�R����:x�6&f��Nim����`�H��*w���qfzj�$�����4|Ћ=ZwD
��g�@�7�7a+[,�IL�wн�K8FU�Th��O�i7�H�[RRBl�����D�w���&��vԽ�}�/\L��X��Xw���VWW�������tn!>�5\���x�ne�+�tJy��36��#<�u��!���ܡ:y���X~���I�J��k�^�4��O��>e�&j��Rh��l�����7�Nf�1�hkk+V��{�>^����Xmip8�J��(I�m�C�V�po ��@4��J����))�����v��Nf���r���kr� ]��	A`�L���@[������4�0v��% H߹�����Ĝ��x�aWp_� @;�.�Ycե���k�$��G��fff��{���w��}+(�rt��R��T���z����>`��X
�������.�� v���!�io�����؝���{�� ���W�^,��(���j�l�	����Q�g}�h&����Z/Š��9�$�6R��w&Q�/���<A"��ܢ��Ø�X��A�حI+Ow:���h��奌L0�_�t���x���K����@&]EC�C��ۮ��|���W[�W0B�<���;3:�W+�j1��|�xlA'����Ǝ��Y����>6ϭl�ߏxb
b DG��:D��L a���EC�ecxyy!j�D8����5��z��H�k7���{��0��^�63�м[���!9�h`�)~�6u�#G�|�;e:y~Φ,�# ��!浵�\�4L0v`> $NC�W����+Q����O�@o8 �w�6�r�A��z���[Oj��Qc�|n���K�N r��R%�k��#55��:{j���6���T����sMD�Q��ќr�[337�ogH����)i�@���0!�����]��I\�@��/А��i��P;I����n�����(`��J9�����D4^SALWxf}&rϻ�� &��?d���'z���b��RxI�7@Y"�J�#���bK���A��̄����'PO��I�}�~�w{ޛ��? �3�i&�l���ˈIJ
��ANr��:W��I135>{�0���3��}�ѓ��'�1^�L�<H<7`%�ݜ��'!$,�2y��p]�A��wEXع�4�$��B���c��:d����2

�4����L ���G��l�x�� ��7@����Y��m���-���gɬ�6����ё?�ni������b-�0P��c�w��r�e��n�CV�eM]]���������0@(g�W�F�	'IC�2���HyE��5��i��X��s��s�՘3%XU>>Ë�k�|�=�nu(k�:�b���eQF�������.X�i��t���,+��Y���H�ä���RN�_��B2���˨FI))++V���/e�m�{5�3\8⎺�ѼJx�V��:p `��6�{�7�G''���w� <����E�.f�/`��®�7iDk�"��������K�or�+�ø�ڒ�2p b�N%�5���]�5XS(?Q�1��;"�}��1*<�ƕـH�)b����V8cӁ�I�- pg~~���o��`�3�%L��hd�[+u�%�{��RxPw��B�0͋􌳣�b�����X*iJ��7�<��Ub@�c���j�R,1#��P��X$&NB2�}E�zDN�Sͯ�όҝ��ר�3�]�^��-2�7��ek���Q@ �*֠!H���J� r��慅��V�ޙ���#բeN
F�����c��l d ��G���ٱZ�zU�����VD�;g��J�^mm&t��+~�/oc���9ܣ���ʊ��ik4��=��Q$���Bϊ>8�� {*!fv؞�����7"����IINF:.9�p7 ���E[X���e��\f�ǫk�+�X,�`��bc I��O��b
W� b0���I�_�����|K�v�A̓߹� ��a�3֔Jͪ�{�Y.2�8�V��E���������W�?땗��,�7^���Ðf�_�=~�ӛ��E�?�\�RK��(\y��⽂�R͌�WT0~��{�������5[�Gi "�F��&O.�ɫ>&D���>Ĩ��t���0Z�x�.Ӕq�_�鴱+++$�,:��5����˴�%��%�����%ask��	5 [�;,8�����f�4{����Sb��KMMO���I��t��UUUDQ��������ͫ.��
�n��t���ϐ/J�^��Ҵ�`��ѝ��x�		]���U��H���^�U]]�tI�wP?oLM�����A�����yDK���	������]%����lcrP�"򬻂���_dfd�� ,,�}�2��{`pK�T/�0�:�����S��{X5ɗ9)u����m)%��_W��c�@���D��h�>�����5`�O�oGG<yp|��U��� .`�J�9r�`��6ݚg� ,�~Ql�C�G��n-on����n7�����������	kt������W�����X�	��������?^$�����j���!���h	��Ǟ�t-rD�`��Xbr��#WMCI)��=�*�?|k�J�v������N��ń��8׆�āZ�q�=:�����Wq'��]H��C�O� ���9�����?baqV�6�Ǫ?���$`c\\��D�)-7��󫪪���5����ɖ�����U܄��T��:���K�٫ey@�죩i�����+&��X��0L̫�z���\0BM2���r1r���~���C�L�H��oG���Ί:�@�����dK��,�b�9�Gt ��~Ħb��L�D���^�W�)1�u3�m����['�*�c���>����9@�:6�uP���ꮜP����1f�+����}��DY��t�y��;~���� #��ʖ�>�w�K��Hlp�'��E��/>$�+1�뽴<���NϬ�4��I|�e1=���m055U�͌C���x^-w�.���G�6�y�J 1-8�Cw�<����s�73.:%�E��i���Е ���>�bA
�F�U0�&_j"���H���+$�
fԻ�ࢇ?�A���eqX-�;=�>"""Ҏ1�	E�����x!�2�Wl;A�T���3��Y����Y�RRRiJ�2��X�r���_1($| �(�:�Aa*�;c���t��$��wF��`Q���g����&������{IOO_���񱙹�&�*(	!qIz-6�N�x�MW�F�V��� �,@߰Ȥ��9��~��u?����}n>>2� �:��a4aEEE�n���R%�݄�Htʶ�����������l�x��0�=�{zZ �5�?� ��x�J������`
u��pε��(49��L �it�8:;�4�&Df�HC�������� =H:o����?��A�A�A������Ջ��p\�13h���[��6~��Hw���ɛ��*_
t�'���*�\��o1b�E��oD�kt&�?������,��$��f�����~�AՄ���[�Ñ��@�!����x�y�����3j�[����� �x@��v(c�Ç�&v=o_j5%�γ4����_7��x�fwĳ���<�ر��L:t��(*R^�	HI4�O+M�f�]�;���<�[q����}^]]]M���]je��}���8�I\���P�t�
�A� ���]��:�OGp���uc]L�f+�it�>Nӛ����,���;A�h�����3u9�ym�A��.Q�M6���1�����X�O}Á�=�� 
���O,�,�$2�8d��.�-�:cG�r5��X
�n`�*��A��2Z�c^�!isY����d90�Y7�aⲴ9Vb�H���<����m9Zw�	n��چx�$Źg;�XF�3Y#�����zJf��i.Y�,���6ǝ`�C�;��=�;]�r�Y͆�ӆ-��ӆ/��vr���%��
�eyL���x�#�����?�o�����l�~�B\�EA�;\��4m9ç������3�#��xaǃ������Q��(*��0�
_!��l�VG���yf,�z�>�M��OO��|�U�����Ȧ�"��	��ϑ�P�4b;W�����*�@����m�ܧ����h|�m��0�]�hNj7�[�Ǟ_�W�[�up؜,|����!#�!US�y^hXS�����oY�(ذ�F
������5_-���\��_�Ӿ�S%�Py� ��O(���w~�b�h+}tĐ�*� ��c_�� �8z.+N��#�9J�vH��b� ݢU��9��*�<��:�g�Ki�|��c3��S�^	@�tn���x u(��ѻ�
�#����ZA�����lVV�\{;����K�E.n>������.�����'���I�s�Vy�����<�ł*�PQG}�4���b������黡P(�@�[�D�S>�SgW]Z)�o|�jK]V�̘cQ�~HM��_�=��$���(���j�rr�79p:l~���y�O=j�i]�=Gf�+�<�q��G"������^����%jQ�RU*��h�V�@�m��P��}���\�����kȭ��'���qI��h|87�'^vp�͠p����~N!E:���/>�Z-��3�I�޼����̳[۵	�,���^�\Y�9>C=�q�19�y�~4{�f�t?� �r��D%�;��R�^C�
깽7z��P��JGvl5�N:P��b����F�\�)2��O�4f<PY�uxא���Ǯuإif�����|Y��f=?�:�=��:�>�GK�z�$��= ���^�����v���T�ǢvD?[�{��'q'�R��ǱGu��;�v���wO�Y��4_�
D��񋯉�L6���y:�佑`-�Ǉ΂����Pc��Os�//K ������X3�2����br��i�7JT���ʮ����Q�m4��W�zJ��ɰ�d
-{d�X�y�����C<�����-��9�C���Oyr;���9������G�f(`�g0�
�èD�`m��S�{5�_��������A��ق7���xeF�d��C��#ɨܕkw3\Z�OO ���t�-)>�tyl+&��r��j���/�s"�M�b�-Q�n�Sђ��7�`;_�����+aS�(�B3����-�v�=�T�w��y�_���%�V7�n�f�YP��Wr����h&uPx�J��W��f�9jNM�B3p��b|t$h�����Ġ��vsd�ZOO���o��-5�>%F�gaQ�Y_�ݏ����-�z�$�Y��[9h��aP��S�1'D��V�����������`�-�%o�[�?L<K�c�ԷH��G,w���j�^�1(2xxc�������H�۰���N:Χ�N��=\�:N�T�4]g߫o�O�m�*|�����$��'꾍EK����j��{�k�P�4�����c�L��+��$l��7��X�9�[C_��1�rBn����>VІ"��r#5��l��,�����k�őb8�zjo=�N�����7Ț�	�+&��g�-g���0oFg�͙�o�@G�/���)���B�٬k�j)|��?��b;%�AϦ��}B�Wd�3�\�zC�po�)�I���v�*tV�`�ҭ�I�+��JˌM�|p��u	.�v�x�1^�x�q�n'ً��ʓ�9��b�~�K�_Y�e�詝�yB	,�^ܔ�D�H ��5�~�ҠZ�8x:�".}y&Nݘ���v�<x���E@G`��I9�@*�%r�-�62eG��^��� CrãX�&�sG�5Q$��P������/�"���]��t�;������]<p�1!!xee%&6�]&]%���oq�s�m�W�|���(W����6<= ��08�Et�(^j����K���4D��2�z�Z.Ym�C���L49,44�u���[T寮�!����f"E�[Ra�!j[�5����p�P�J�!�S�`߮`@�ڜ+����Ȟ�&�(j�\��G���-}�D�m�x\U���XR������ߙ��Vf$��ը�3X�g�\l
 �����?t��y}�`�܌�a�"��+T2� ?m�m�&BH�=�����A�/�A3Tq����$�,aR���C�988H����M.������hzW��/{p�ٹ|�ܼ�� �X�Q�7��Rh��j6�N�9 65넜I��F������ەEl���Ԣzgh�޴����P3�oj��˲x�+������
	�v��eG&߃E��>�X��L�u�0>���̹b�\��9���N9+N������^ʜ�g�w�9����i$���LGNN�)��t2�u3++V��%H��J��`D����1��	O�~����5Cj1�������1�1��O6�;-���4�ɨ��V��]��}w��w��		]OU�d���6e¡�k<B.u�L���Q�(���@��Plա�+�cG�'��5��̈́�}��3��ML����#�(:nm3z�w�C���Utב��Q�����}�&�}���v8Q�%}���:,�f��'y�����t�33�,/�v�λ���F�ݒP'H���'z��6������&����2b��
h���S�~�Or��w���۝鲪?9��icn���Bso���|�G)/5����.+A󷽴&?�l�F���El����U���|���t݋�o����}�s��W�.U���?~�N���Q�l�A��3�26�n_/y=���m�a������$p�s�8�[���v&7� )֘
T��V-}�.q�so�4�7�<�vf��:�x W�&�D����S|������ݔ�T��PEh`ɖ�)�a߲k���Q��k�W�igTz�QGG�q��g����<�j�ڴ9�����w��1l�=�*��*]�A&s/�R=%��{���n,���|Btj�����H/�a���+�����d!�0���{���8�Kd�c����xu���LE=�\I���?��_mX�9M;b.�0�C;�B�O_>��&�ո����iN'�"1r8R�@{�BV��O1{�N���Դ�qe@���43!���h�ߍ8��'`�4��Ia��P�X��9o����]����d�4{zm��X�r�h]���:=�:w��*9+S�?�D���Za�s��hE�F �ڑ�߾-������,,,<��<n���(;g.d��Tw�]//��u��,0�W̡��jJq�#�|9�\�R֥ n"�&���:�:��H��޴��N@�I����m0����$-��v���*o�##�`�����}\�㝩8� �[3u�w�iĹ�P�|�b���t[��p�o}���A��Ь�B��j�:�d����p��l�AYN��رw��u�Va�O�X
��ɉհ^8�M�4===��� �=1����s�=����e.ך_G8k�)}���sa��A����کZ���j�bՔ�lf0�Wҋ��˾p�F�J�=��YVV60?�(i�ܨ�z\�|�����x tiIËɻ��>9c��+�.����o���v�q���'\�O�F���������ZuAD�Ύ�
�`u~f���%��zb��8W�EV$�*F%5%b1�9s.�C��_�e!���Uh�̕o��t�1�t���mz�~,�P��_j���6������o߾}H��n	$a1>������5��W��h
��)� Q��-�U�wƏV��s�c�޴��7�1LQ�G[%�be_�W
��Y~�T~ʩC���'\�%|��p�2���Mz�xH���IE�0��J�8tbb���E��<��稨��r�����׾k䐔�딼���Γ�����)1�����������3x{/�ίO�(�4[�o<Z�M.�����p���vI	N닅��?w��VW>��S}�˨�>�e�����<�j�~3����o}���;5m$�*��f����jӑFԒa�o�AO�ddd��L��`������> ���hN��NB�y��t�Um�#禮��<�4@a{���7S��͡��䩙!�����T�j�)5b��7�Җ�w͖��l3�����>�n���Zu9mFy9�4!�}�.yf�����xI,K̈(�#������R
u_�ٵ�ص{G?�Q��V�*5���F�O�[P޵�4P1�7����~���@�T�eO� ��Yr��k���$x�G*����V���h�w��ɤ�S�pss�2n��?���ה��D��j�|��m�TLm��V�������/w{�S���U�).�#�{dR��w�*��z���`ϫ�
���ȷ��y��tZ�^��07�ʚP��_%68r�1U2�LqS�D
���+l�ˣ�V�ǋE�#�Rvvvf����8��׶ƀ;ji��Y�(��D�h��֭șMϑ�ӣ��u��;��,��YAM������=D��aV���5$-N��d��X�_ Ap@.Q�r�<��t�_�a~wL�ڠ��ڗ��L��ƈ�zFZ�uU���JJ�G��[�3.ޭ���[�}Y�9�0f��k9I�h�Pl�>L"I��=0��u��򲲁���A��a�G���, �,Wy�wL̚�)�k��#�Pu߹�/�1׿:�[,U1����ᘵ�?�2��������U����L#M.��Y����F`|�S8�g7WM�C Y�e����/�e��:�����&[���ْ��7.�7S�1���w���gGn���x����
���7�G�R܍Wh=�n�aY�[�Ύˮ�ig�gPD���]0`Z���쯹��$'����q�#���,�>����y����fz\_�M���0oKå����_�_���H炵)��;31�$bo}�@p/us�'�ٍ�V���4��m ӧѰ`C��Q����:}�pA�E��
ջi��?�(�t͓����mB#�E��7J�TN�<����z�ӧ/^�X����Z�:Jg�1�0�t��W�0#�{�x�5i988�kT�sH�F'�Q���:�Q���g�.M�Z * ��m��aA�u��Լ\�i��,����
��g+�ʪ�%_~�\:9��æ\��\��)���@�i����[�{�T��v'b���J}2^6���yS�z5��?+hB�DH��F.^>����T�G�P��v�k�k�f��L�3'���y�Ji��6v�ߍtP���������Vpp�������Ƙ���������Ns8;�!�jq�@�K�-k^�u�H-l��h餁��n��@�;��L���W�=�&��H�m����E�,ɰ�c��m��0)���P����=�N�����R��5��� *��@n�ܓK�tJ�YX(�%�`�q(ii��yK7�b�6	��<\�޽3p��׸ɶ<�����)O
�n��\mϙ3�9ў�%&<?�,�}2����.��s9r�z�r��|	A�Mc+&�YU�y|��)����sG?[F�߇Ey3L���n��n�$�?Ǥ��^Ƌi��"��@�G�j��gbc���3˷����M������W5 �����R�Kn���J���"�55���r�[���a�O���q�"�:n+U��쳟�l��X������,���ep�a!:Z��I��Q�3R�U�-���w�Vg�8�ޫi1�`;������;��,C?��`����9��doc�jh���d��n|��{`~~~ ;89؈��~�b�  �҃���@���q����<7����.�~��w���5��?������e=yW.^������d=�\��U��p�~w.P"��׹E2����݊y;D�o���<>����Q��ٸ�w��߃
E��oVO�z�Q�Ɔ���y�p���k-)�*�%p����XXXT�1�%%��_ F���"�)�V�TMz�	�+�<������q���ʕ��{~��J����0j~Qgi}��印	N�OַW(t�@��h$ҿ��@5�U��T>��&l���:ɽ����$]� �⛘4�3Z"��̯����:��q���� ��<V�_N����VW�����o����/ ��}�G��ӭ��D6A���$���:	Ȇ�"��@��~qP'�}�V�:Gr����HCPBg���p%�A2���k'h��V!�ע�=�W��z�^��
d�x�U���N'Y����A��T'�&���n�6pc6;�ef*]N�ɑ���y�,'q6�H8[�WI�vP��O�̱�'Yb�1�
QWW��a1p_InP`������	,ؐ�<0o.k#ygA����bnKCX���WI���M$Eկ��#G��&�K��)�P+\�S�[W.MnL1h؏9�,�G+��Bv%�,؎�l[�-Rc��oTx���֖K!e��x��I��YII��y ����pm��0���e��'1� a[��ɂ��N��P�T�z<�]եf���]�6������G�$�/9�:X��w>�`U�$�f�fJᑹȠ���+�n��"�o��਩�����y$�RX����s���D�3kpa
j�|M�IP;�a�~m97m�OS˩��=>2��q6�0�o4v%�M������x�y��O������]ӧ��rԦ+�:9\����VIp\�F,�z�M@�¢v_��Uh$�)�;�[Z��>����$�+�.[�!�"W�l+w����Ĺ��Vt賑�OSx���U��M'�dCդd�[0���%钣3T��Zs"��5[�7a��^>v����4�S%zp���e�A�DO�OFa�ͩDPR|bRR��"e�ɋ�Q���f~ �>}�$g��zC육;��dPo�|y�GO�9���E�7B��m��^ý<��CP/FC�/y���j� '���C`3��ө�ʹ�,�C���]�&s�Ž�I��`5�*��Z����b��O'���ܜ�M���4mL�RR\\<g��k#dm�)1��\>��}u�Wҷs� s�6�˚����l��'��{�8�nŇ<���P�+ݟ)�����e{���1�+;����P�(��v�8�A��$����V^�	q]*���H�㞈�q�$k�\��9�C{�P¢�=j�:���i���N�V���e���v��ݠ ���%��+:w�)�L-�䔙[���|��3;;��y��G}Ν�F�/V$c��%1�f��e��tG���� �$r�c���'|T�{��5���'J��X�c���DvW��gټɽ	����,)�������9-D�q���! �� �|��j&F3�S�*�c����nߐ������c���W:�:~Ts�I�P��������}9��M��n)+��r�v�{[�0���B�DS���8G�
�C�,X���"���$�z������<)2:~�ݺ
&7s£��0!���t�nnn�jj��|����Ȍ`�ۂ���-� 8�J˘A$&�x� f��r>{���A�-q6���^���97S /���Y/�Kh�vv/Dx'A����=e��Z=c�<YXr�}~�[���h��k僴ݹ�R�(��HlȺ���Z���f/�S�^��^`\S�>�]��`iOFF&���0��FC�,�shԑ?CEl���#[i��g���g�Hg�+y���Z�x9/{n���=�?�m���TYe!A�'9�A�:G�.���kڗ<��=�0>�Y)Z��kCt��T7E����~/���hƂ�h��Γ���+���o�R�y	�/�����М���2�բE�Shvv�V]���+z�����d� ۔>Hj�h�Q��/*��-q������ǿI�ߠ���c����WG`���.\��bn�|5�H��C�Ǐ����W�mz�Ճ?���`M���]�)�R^k�*��6��a��Ͻ�3�^��<v]@�����Q����SN�G"M���B�nӑQ���� ��#�sFdZ;- �Q�y�����6�b�F�\�?B%�C� �Hy`a�ڦj��Myw�s(er��r#	�M.[{�oU7D�#<%�%�C��IfXÌ�ע�^�{�cK���Λլ�bG;Ͻ��$F�%�CF������G�ͫg�F�Cn����w���X�7����O�i�v�%P�6=I���a�tci��Eqo��yLN7��^\+?�y�Ϊ�H�Ѭ�~Y�8BVi��?wZ�c��dS��T�B~>�]�-�OC�gg0�{�t\,>���<�%�Q$��)�=����98��n��[n��o��mc����w�9�kl��Y��w���qzP��8W�:�	|���B 8��l�������)�85�M�2��+ɦ�z�W"���Z��>ϱ̞����47��)�Y�jk�qgt>��cwSc2ԧ|#���= ���ә�X7���}+O���c�S�8>>��TL.��ڨ4��m��<�
��&�,��Na۸;Z4p��������MF��[坭��YFԚhf�%@�J�u��:�΀�\�|�c�c�n丠$YU�e3_Q5*;A��5����ι_�0��b�2��K��{\�n����0$,A�����������DI�(�C1ܪ܊PQH����?IC5���������ڏ��:+[Q.�ν�hfy��Y%d��?S��5���j� 	R��7���M�~��&{��Y�,@��q�!���A���J��2w׃��6%���(nHN�d=P�y�__����V��\��f@VIf�U��2��o.�L���d����
7���ּ-�}J��d�}p�c�E���z�63X��:�Ӧ��~3���������D���pYP�������[AR*S�%����%��D�rKM�:k�?ܛ?��O�7j�[^���;��Z^Pn6b@q.MH1pI�5��ȸ��n��f��a���3�QI��Q��%�e
0р�?}X%+#���B�c����IЄ�B�+��Y$P��� ��4F�m,��>R2.�����O2h��4����i�LQ)^�f=�wL6�����fD)GJdw����9z|�6Eml�2Iy�����dqs�����3'������E�A���p���>�z�D.�\�T\L�?_�P�x���H��ڝn���o|dh$��7����QN� �{Ѷ�i��z�B��21�[V]�ثfI��n�ދ9��=�-Ā�)���x� Bt��"�?��Rz����ƓS�2x߇�T�K�������a�ׯ_L`��-���+�B,���~0�ٯ���a@�v�{�'�\g$���ڟx���#f1Y�;��N��0CFL�XX� ���� +U����ء��9`1�yh\u���\�fG>�\�%�3��c�=.�̬������-1�ߥ�G���ߎXH��G���b�r�t���E'�5 �7�ؤ���DF�sY�V��ܗ�w���L��ȃ�j�>Alll��ǹ;:;uK��r4�e�U�wF#��o�����������-i�m2�nM��4��!���:��yO�}��VmD@:OMX�bf�m�_i����������)��n=�Zd5���Z��ͥ�ٯ�����C*JY[[���A.�LY�:%o�*v3���g'��X�Cu�졀�d�^�2��9�m������ �܌��zO�M���A�ק^���϶g��R9��3�I�CBB�Wnfɦ��U�{�
8�6%NDmO{�E^^�Ł�T���y�N��Q7Xb�H�d���@�π�thD���^�N?@7�M��)g���J��<��Q[kB@�[Ȟ\���H�q�L�;�>V9�F�&�B��	�f�b[���t|p�ȅ&�ѥ�\��b�}���:qXj9=��=��K�]�ف������k`�}��`�"�hx@]�b�Wh7�h}�&Mdp�	I#W���{Iޤ�Yg�A�j��F�$L��q�n�d���\6:	[	�D�8��i7}��+�9\���?#��A����ϝv�Q}��V���:��� U �u��0
O!'�->B4�5߭���ț��n{e�j�:H�-Ԏ��7Z�j�$j5�3�Q� �S<��XF3���c&��b��$��B��I�b�x�5��1� �V@4%W��O7��D��/�� ��nlD2*���)))�
B�G���9��T.V�vvwa������V#(Wf&�~�b祓��CC�HkN⺴�b���h�5�� n�"�!��ݑ����45!�Ak7a� �hɅu�`�-�*k�/������C�M�D�OwFs����>b|��2�E���dx������u�+�Rq/u�MS�_�����1���Z+��-���n.�<��0�X�@�����1�}���C��TJ�����b�Q�+k��1�=�FH��vn�5n��D�'������PRS�@|׷`DYYٜI��׷ЉP�e���������[�!5aa΢L'{�܍M�_H��.n�1���^���T @��7��uٓ�ho@�|:�.S�G��f4���[�|uCMe����������V�l�վ���>B���hSsyՙ��ׯ= K8AQl��,I�����&��m�ɼ���~��n��l�^��B~�[vF6n���Y��a2���2��gגo�4��N���T�쑻�:�ݚ{hҊ�B���\I���8�C�u��Ό+���-�Q��M�Ca>0�W�/#�t	�yF��z+�����r���w�?��Y��SÖ���.5��}Y�@ؑ��I��{i�ƪ^r
C��yxxh�X�]��	�\%���"�l�k��E ��Ξ���!Gr�:�
����0�|磹�HK��U����$���>l���ޝ2�o��w'���b^2T�b������ߋ���\�1^���9�$���ȏ:\j�\'}��Y��4j �2����ď�b�� ,����l�e$�U��0^&��˃�l���g5����l;�j=�����0��x��vܧ3��(�h�������Wx��Ux�`V`~������f�%?H�\4�;��f�2��w�hZr�l���_��7p���)��S��<?�濥�G��Q�(��:oC�a5�Nz>>�T$�4N^�[�ͪK�$��2�\�q��$�]~����2ԫ�����ͻfC՛���z�e����dm�>�>�~h�!�FaLtc�L�s�{_\}?,��j�[��]�Ƶ�M�=	�6���b�L؍]>$I,K�
7���TPPHui����n_i��O����� �P}��7��c�m6�z搂+�=11*�)��B6����zpd�=�`n�a����#�f/��ET��py��7iڽ�#Lq:H�=^��T{յK#JSVV֭3Hw�|.?[#��WwEJv��������믣4�M�[��]���z@̛���K:c$����#Jh�Lh({���x�����1�6��/̖�i��H��
�@.l�&�>�ɳo(<ǧ�<k6���:�B��w]�,��,̞ɵZɵ���fQ�U��]�f�gǓ �Ϣ�`	Ȳ�����:Ma�	��)���>LhB@���I�Ď3(�W��x����'��KO6�+��Fw��z�,���QJ	�g��q���Ϛi��N�N�&�kG��s�>\���y'e]]]�G5ݰSj;x%Ҹ�׍��C�$����D�K� Ɩױ���BdQs�n��������({Y�4Brn�r�S�H�7@�������2�5�������4�v�aA$9�C�s>q;�&�s	"=o�o�����'Ot.��S~����5k�T�R0�zHL����T�K.n�@������ ,x����r]�b
%L=wP�\�������Rv�P1����	v��\,�aȲD�����~i�|i�5M;���l��{�3� ��c�
���`ێX홿;2n��ܶ)6����>��\ZXh�!5MH���k��o7��C�g_�EZAZOBDK�0�X!��ɪo�jܪY��%�F[[��*�'������hhhdhrt�\��%,��������n�ø�
���m��������|� ��/W��w�,�I����1<=������0���S�**�Wt��|b��W�/�&k)�&�OĎ{��燒���*"��c��|��*�7%A��D������_��~f��
�u���e�^������q�_S�u��и�}6�<�Q�7 ���<�L���w���5V���{��Sƃ��֛��X{�&�>~�>�PZABD�.EJF	H�� �9�Y()�!�膑<8���1@Fw7�.<��O�C��u�5�}��O�{�]}F�3@�8L���ѭ.�R�;�����ſ��>�
z4$r���(#��Ed����D?_Ƚ�9�jנ���k]��
``�=��4�>� ah:�(�ӻ{#84�kZ����5`��Qm�y}V��R5���^sV��&B���\�~z"��G�@�
��5%B!�Q���LMO"Qn����B�y�����K��TR��>�C�E`ǉض��-2XY����D��b�����Z��8�$�[z��_�g�E��^��[X`_s�# ���4�f��X&n~��~}M��GBǎM��ԭ���_X�R)����HN)�iWN�E�L���`�"����5�2�jiP�(ŕ���c��� ��DG˝��Ua78"ڇY������e!���ƽR7t��
���� Fqg�T���k�L���+d 5��D�d�x�z�Dy}�S�:��6P�]Es#�Uyj��x�R��1\0��mX�ѝwN����5ʖ�f6�4����������2
�6�rX;az���������	/�:�R��iػWF���t|����e���"���dffU� ��}N�]�jf�*1��RG]ȳ�{�'��oڰ�)Q: �n$x�+��Yٴ��ne	L:$��/V�샟�����g֏������=M�����d}5޸�jY08������9�'P���-9l7�.K��w���0%y� ~���u�2��F����*z�H}(��d����C��886����G�X����JYg��D657wљ�2��#!*,��DK?/�Ժ�ùƋg�`	�3"��؍�Q��Uf���V�+��ʚr�1��ݡp0��ӗ�c�L�FT�9ҟ��%�,����y9���C/�u6��žEŷ_�xv�?���y߾�A9�i��Ωq,����n�v�Gk���D����	�����׻��]�6����R�cVTU����O4r+�9V����P!�ߏ[7���Fó�n�}�S�-��"�R-��:):�((*�Q=�" �aV�U��ܲT��A;XZu�ʹ��w��$8�^Ç�_5TU�?�<�0�^5���l4U��G����/.֏=<�]s8��D'�8Ȃ�W�^J4����4�{ϗ��O��w#�jN3S�q��]�U�P���A��\�OP�����%�CE�]�+�fK㻽�Q@�#*�L�GO?&(כ�{�dSH��	l8=8���ܕ"#c�"ݐ�t�`�Р��YB�g�����%��1��'�~�Dm�x+���>����@e��6��j���*���Ǚ晽]�y� �
�.'��M �ڴ*{舘{��~�����lhR�މ�S�KJjʆ>i����`F ���/l����$�����F��l����	n��i�m�+RBBT���~ݥ�.��+#�!%i��q"W�/�hw��S(��.��;l����7����!�LP��]�"K�:XȾ������`�R��#�t\	��;Q�6���T�r�>e{�҄����6;���:�ГNA�-��״�;�z$ŷ�BVy��eD�4�Ud�7����X��Q���V��:g�l+J�4���V�������/� ֎�Q���������<ƅ��/���Z���*��@fy0��������&E	�����Ŀ�뎶QD2�x�sD�3��]����4�O�t��X3�d���yN�EG^d�є��.��_Xx�Ӳ��6�ܲB�u�[�[h#$.������O�y숢���P�ylA�C�ŉ���Y��`���GB���4 z�[�l��5�J5�5�����e��+*�,�r��'��ݟ�*�ߍ��/�O�'o�������<A����_H}\ڿ�|��~gR���/�����#UU�`h�1�@S�p>v������j�=�E��ϳ��Tv��m}xL�ĹΤD�.���_��u`j�$���
�܅��1Q0A����*XH���J��l	�r��"՞h���]���w#(o���t4�1_��Ǵq�Y�L�ooN�(
3�� ��|����F�%���Ja�R^��_�*���*�Y��a�|�9y��4�+����`�ʏ��ꥭ�Jqk��o�/V�)i�����`r����y�qE�>M70k*b��;������k���4_��s|d&\�_3��Z0�Q=_�c�);$��)����$#Ż,���;����
���1O%E$��ՏP�8��{\�;��t>�0S�3]RL�Ϝ����R�C�U�������#c,�j���*�>>�ԅ�|���*�7�cf�ӻ0�6�������}�@b��x�����B���'�3���j�W;T[�*�ei�f�[�-�\:�	Q`~ˏXsy�����!�D?��bL9fjK���=�('�\�7|Ǌ�&\NoSk�	�y�k�r�n�Jr���\l_�F�È�2:XW��G��dL��`�q{�J;��:S8�>\`��Zы6�%��;�݌.N�NxcU����J~���C[���-K�;*v*v��ļ{��MZ��!�Ġ��X^V��Z��<뽬o���ݫ��\'=��ȯ���ϗe�,Wu��*!v�12��w�>���kI���z^��M`ۿ?�(ﷴ^E�Y�D���|ޅ����ҵ/D�:�U�}wiX%jv!q?Ȏ���c�������R�!���\n[�[�ֻ)�c_�Z,h,��Ϭ���G�|��v�\�V��^-6����IE�Zl~ܝ���r[��i���=N�Hr���u�^��
�;����|hy�\�/������oa�m��C�+}i8'.	��R�A�Jje�(R�mE:��w� �R�o���콺)�����$���:T5�\�xq;���\�/˽�������#��-��f�RWFE��z̽q�Z[�����e@������3�&��O���ߧ�Ȯ,"X�\��m�<�:�-� 5��<��X��������M�.7x,Di���{.9yM�_�A4����0�=��
���w�Wun���)�
6v?%�Žu��}��<����+�2��R�=&�6�&�yǾ���_�Ҥ�3��ZA�U[��]Ǹ� SI�/bo�{�f����}��n�)�eޫ_&��d�Z-��{^;Z#MW��^v`\:E��q��Ҭ�]�O_�z�Fʗ����C3W ��?1�w���b��`�lmm�,[� M1�ʘ����d��;^�)ι���W{\��В�ZֹN�w5 ˹Wu#W� �N���D�)S� ꭏ�SZ�zM�ձ~���I����&����6s0��w�e�����*�bC�m5��b��ư���[OU�u�1H���|5�Y��&�<��w���ݴ<�8r�z���ȬRiR	��ڵ�m}e�c��7h �B6nΠ^��kdTϋ�8�.��}�nâ��ūdWCxQ��O-���e�֜M�8��@���
����D(w<=x�ܖnO�9P�M.����_'X��-����� ����6ɑ[t+��W��ڼϲ��ձ���:n	��yONa�_+��s��<�oXr����$�{q�5~��S�^��|)J��z�a���v�[b%���/��w�X#D�ww��e�Hz��3���i�3�T�*f{�p�{ؒ;�J�ɖ���S�	�e�E���ݚ��6�H�V�W���y���*��<Bz?;`��uQ
jO�(�̶HNOg+�	����vU���xzj ��f'�l�z�U`T��?\$
n-RG?p�w7�@P���ӽq'5�!l��%�}�����.�eoh�H=��Q�d*�)5�K�s�օ~))����8l�4�E��DjۯY���F9Cj��������Y�eBN�;�mAJC����4���lL���k�]0F��T8B��{ug���{��Z�xz��	lt�U��^��_L�0\­i��e!�#�	5L��ɕ��ɩ=�򾐱���.��k^��Ag9 1��\e2Q~PZY�}�5b��22�s�i�u�>gN@Ί}W���i����c4d륓����ܖ�Z�Ӧ4?���ͻ��h���� WP���\�g�'��bF���׊
9��%�}��_rKoO��H���C��S0�Wr�E�m�`zC����ȍ9H-��L�x��t��u6<�1���\�W7|D�Z�ؔj_:<�9��@g�q �O&ظC�v��N�g]��IQ3�]�}1������ �8��h������e�(Q�f �"g������*i̘��o��R�Klv��z���Ĺ�i6ƹ3s�Ub��#Ϸf����\�q�ON8��
7�L��u'vq��5����Xr�F�7]~C<����!MeE�Xu���W����s���X�k���P���̺D{+��]�l�s��3�{�5�%&d�/n�)�C�G�4S��6	W�XYl0��ؽoSVZ���ӉY�В�w3' !!� ڃ��"�m�Ҁ�iv�*!����nwJĢ�\l\��o�:�oM�C���B|�������>�;��Vh���[d:��#_� �2��¢�����>D���*��B666?uu>ʔ_4���+Ί~����Ƌ�L������>����.(r|��χ�<����nT�KI�f�B��kN>8���%�}�oX�X�-h�s��PH�c&H��9�ɦ�ֺ^����d��`���9Iv�������U�td~��<�s����xN��gV�N�g�tR��\�F�I�XCi�ֳ��\��Ҧ�|�%~���<���#�u^���dI�]��NXC��|Z;��4�j����-���������?;�w������y��$�n���<-ۆ���m�K����o�2�������&�mXh��K����`6 c�u�!a��S6'~�P�?$���O�; ���P�~i�u�	��� �	 {���uJ����
�ů|dadcQ����>��>��;�K�oh\Yt�RbωB�j�O7�p])�|�u���q��~�v^�MъF� ��R����N4d.A�i��\�r�ٍ.���ƅCM�M��ǣ�X���v���~o����76#�NVVV��D��7�`cd3�^mыo߆�ЇIii��n����_�Srr�"�EFN���'� �B�233�n�L��	No�����\{~�h<��ǯ�t�Kߟ�r��S�eD�h����r	S�0�wk�?Rn|����Af��p�Puvv����\���			I�����������k5X�Gf�����bT�}�E�������$��%}�� =G��(�U��RZ�x���P�x�9�r�=K �m%�� �P��F48ajjj{S�___�����C�q��V���!<���-п`�1�������O��O�	����k��}�$�����̬,�r�E??��z�#3~P0;ê�'J�d	�}7yn�S#��y}/����ఞx��@���e�e�j�����0��R�uQN������=��h�x���jC�h^f-!���#�'�����f*d�a�==�-{�@CW�(�kw�I��	�Dvtw�	�ek���G�.��`)�MO�6����5@��n1�Cc%l�H���g3[BFF�.��C�JS����������Oxv���Cg�\��~�N�S��5q}���T��o�{{������X�yM!�|�6�`S��� !�2�ܘ2��������%Y1ɝ���;al�sU�W:1Z�M ���Ȃ�s��2���}G˥+���N�X�9�=�L(��.,.���r��=z}55r�ʅ_�0F3K����UU���G�z���ҿ��sC���(���i�MO�g��g�-�(Aϋ����kb�����K5�n����I��s5I��㎉�u���F���BX��XH�2rsoG����1�� ��)9�I��5Pꦺ�����ϖ�\r5�K{�Cn�}_�q��m�2:}�{�i�a3Op����kV��4ӖD����&L�sssk����K�<��˺p���T��v?�i9J�:����z���])U{�Uʘ����k�^S�ȵL����oh�����J����H�a����'� e��q�a0t:��x��h3�����i#�1z�"=��*
��p0�Ȏc��u���u���պ��?.u�,aE�r��Viq�x�iyR��-?��W�D}zj����+�&[��R�f	�v�λ�Ɋh'��<^��+%�bƳ���u��������<�l���R��3��}Y��O����Vƪ"��.OF���)�Z�����-w�<��`�?>��-��a��赝f�Z���':d��w��5�Fэ6�f��PNg��Ǐ_
/�=88h�6�����Eƻ�3��.����Ф��	��#�C����{y��US����4SH���k�WV�a����9*��G���e�m֓)�Z���+�Co	�6Ο���Hz(�q ż�]j�<�_��0���Њ�w����T��T�v�����|x���5��vw���wc�F���	,�B����l�RSSUTT�I�e^ ���@r�`:V�V<�~O�8Y�
�v8�pdA��o��Mg����D��n��sm|z�CJU��ZZ���(�nM�4Z�Ga�a��S���KY�����$j@e}�޽��{��.U&w�� U�u�d
�Α�����?8���զ��6�'
�s���:�?�J�~7h۪���8���yy���ٲ�O)Y�%6
p.��s;��y7I�ܮ�><(��ގ�~�%��RǱ�X뫴֒�M�@����{}�|G3'w�lߓ�S��c�`�	�c[�w7����<p�s��G�%�����h���,�, m_0��� (t��wo��K;��a�~�ﴈ\3��� STQl]� _s���&�u�6�0�r������f��`�`gL�wu�9�%,v8�-��K&�k��x/}��܃�7���%������4�O`JOP�O��/''�������(fP��r555�!B@P�2z�aJ����v~��z9Y� ��F|�w'f�����Y�)v�[l뜤�3}�Q��k�8�cq;>8:b���%~���	���- �I�`u���Ut�\2��f�`l�77�Z�:��� 2�	?�;n'���'gd���j��dDCLdl�{%ld��q�l� ��C0vvE6i���:5�ƾ����t�w�m.v���2��֝:_����fh$P�+ic_[0�s6P9Ԝ~d��U����)��3�E�QF�3���B��y���w:S�K�����(Q�M۴oY���k��F�|�(��@SR��?\;j���T�խ�d�q�(Zھ��oj!S�!I�܃g!}����ԥ�7�hR���d�P���H�L�"YR��|8������F=��H2�[;����O�l�o7�|����e��7�2�
x��}F	��ƺO))`�GV�26~P*i�?r��R��b_��w�nf�ź�+*�	IT*V+);�VH~����J�"�%�����6<�(�^B��� =��+�e�J>�n t�E��1f::�^VN��m��.T�S˟RT��u
�d��~��%�2;��˙�EU���C c�^�B��OKk�Έ�-�nD���φ��c�!�� _��~Ei,�[����۬)�D �^m�ڛ�Ӱ!�imO����PUUuQ��DaxrW����g��!}��2������ӾѴK)`�Qɰq��[��e�l�_�C�[���#�뵾�|��0�+C��t����e������O�ҒӚ���|��n��U�o�Fmق)<z������_����#8���6�U��sW�,J�׾R7�[c*��EFDHKII��|S��h*w0n�TQW�@�Pn����^3�������[X;LMt+���J��G`�8t-ޙ��H��6���X�r��zlqd)�͏���R;�_�3��qX0"kE��j��������g�D;��AF�k�tE��>2���[@[�WO��J��������;���#��<%%%� ���ŕY�89���4���7
!$D��d�$�?Et��+�Sʵ�n#LK�@�b�E/�u�����IJ�j|�I�ʍn�hH�6E5s������8W��X#������ONd�V�aZ�lO�-*)g�U��qa�%��E�������&�f���~%�'�A�J�Ya�d�w�[�+���n߂%$$���l�7���N���̬�q���y�\�e�58'6IX�ch2��-�g�:'�Y�<����x���s�ba����,`�Tյ�.�5s|�!Xb%�7�@�Ψ�+䐥mS5�Zx����Jj(Vd�SY^	}6�h8�I�-�����P{�5�y�?���}�Ǌx���qUG�LI�6�귳6%��y�	�Q$�J�j�Avdx����������@M������^���M���V4�J���F�bn�J��-YN�-��Sw
A�ʳ3�2�����g��cP
�F�R�j;;��i22�=}�ѷt�����Nn�����/��x���(.$FG| �����{`�t��u�,�ѭ�%����q�ߊ ��(��M�� �R�EK���u�=@�)G���_3'<}VEB���Gp��Ë�ss�z�مZ�(��l�[�KRb�Ѓ=1UM�M�2�/"���v>�X�tmnj�1ٓa%əP��PPfb��)�_���F�	�輦V�7��>H�6�\�W��#n}x���m���3�#���4���*�3I���C8�#���!���v��)�=@!��"�"�[�!y�9d%�����w�����pO��e�f�P9�������.R���Ǹ7��N����װV�-5w�ƪ�V��@�U\K�Kt�J�9Y�yGz�2Z������;׍��j���2������Cev���`/���;T̪::4===����΂� ��q03��6^�~�z�'F��o�ߪ�w
 :eۄpJKEI9;�����ܓ\g��͐�����%bqcf��Ol5WE��6޾Z������AŞ�J�CuX_Iq��@-G���z?3����|��?�����n`�>�>4���m��y���o�GL�[y�� ȫ�.�� ��Ʒf@�=�� ��N_�]�[%nrb�l�Xw}�s^U�b�x/ſ"�󵸛��� ��Ȧ�g�)n`�l�J~�b�׵|b���Y��q_U��r*��sn�b6�CӒA&��t0��`8PY�=�2��L��t�U?��b�wБ�18#ܗ�[	�hՅ�C����L�W&��,� 17�[�I�Η�����*G� �t/:�E�A��׬�qʶ�l�D�6��Z�3;J���U�ϓq�����tRa՝Y����)@�+���%�]M	����@��W��a0Qrm��:���8`�d���285 �o�V8́V�����)_,��\��PuF�L����F�Ws�i���Rnex��x�\�P�7��@�2�B�� ���>d�w�TX��~ĂK":�5n(���^�i9{=���!2�F\s�u���u=�Jѕ�����=ΑfQ��_&mJ�����Ф=*�"6��vޛ~s����GR��(z1e-�W��G�e��f�B��G�G�3]i���Sm~����B�bll\\Z:�6.DffmX]]�S�"avdT}�t��������V�g�tG.	�sZEZ�VXn��6*���D<���8?0��7M��,a���ћ�f��v��{��끨�;�V�4���mjS���l���4S�
��j�-��]���4���p�D�Bf�*�a
�6�h��=1�16� ��:��)4��tDh���n�T����G|y;�葼���-���ᄚ���ƀ1Ͳ,$Qr��!lFĂI��k˨���mll�Y(��QPP���]�}���;��0C��
�0��#r&�7����F�'7�j���z�R��x���0�
��c�*�6�Y�{��2���/vI�D��-��p��KZ$���QE��!�Z��I�is��;�����K���5�9�< ��8Mؙ��|r�0���)
咀��H�f��o�U����G�����"�ȁ��Q�� �xN����#` 1�Pw﵂Ø�X�������C��ylT�Ճ�ZI��}�C�}-�o�c~�8���/��9��O��4�<�ߧ�6<!K�ħ��d6�p�-��z�+�m�ۮ��O��8���U׏2�`\�]�jOL|LظN���Okkk���&�����H�'���� ]�ܤ<,g� V*����Ӌ'�(�:��ܱ�T�c��ۇ[`��v��P������}䷆��mz�ЃI�+�;��2^�������xψm�*�3#6,9��%tҔ�����Q����������E�j��DC�h�mQ1��5q�����������R*a0"�Ԝl��@�ƹ!&��������z� A�A�Ȥ�x�&��{�#�C���65�G�e][�wdU+��J{�
�0�8+���Pc�w�AO΋e�^���~�[�������C����K/��*
%��n�l���Ym|��yM��[n�������b{�{̨���횥���N�3�rԇG�t���&�� ��o��?iY�-��)*�t�)Ƌ��9߭��;�c�{�A�z�#��a�����'�q�sg?>^'V�L�	����рiȪ9���
��-!��`��0���h�)�"�EH^��X�@�QQQ!��ySs��.D�u��6zg`xްrV�e��')��+�b�i��@q�5�� ����ݻk�n�7ֆV%m���|U����9�<|"�ೳ\��(�JCá]wk�<݈����);����H`�\������4x� �Ot~���Π�ړ�z;2��Fo��U��ڪ�i�<�w#c�+�%e[l��k�����]��ŝ
-�*����H�H������y���U�$ٗ�\��\`�%��?�,8#7���3�N�����𕷍���eA�� ��F�Yn�\�t�b�[C��~ޣKgB�ɺ�FGq�e���*��J�w���j�N�>g�������i)�����\R/и���k����r36|7ц��λ�����5�"�t��+c0 �eeeU�2z�:/Ϧ��������Ѵ��&���_x��{{z����/�}&5��E!��@����r��&���g�}q�ʵ=���S��S����H��n>�u���"�#��7�0� �u��WF����U�.\C����62�5�^��9z9*�+8����rF_f�Ɛn�Â�p$RT[G����t ��������c���������s������IoN������#ԤLG�� �263��'��@by�/���4��=�����{��Նn�Ud���+**����?^�z�z�:��nC�[7����(�I�ɷp�qY�<H���t����=��(mT�01�c���b.��ѽ��/����8T�\������D@�;�G������ 2MO�F��/�����75uu);;;��EYe�> ;{;g�J���n�"�P�R&�&j	�V��U����-�k�q����Jݑ�u�ʡJ<��oG�c�_���@�I�K��͡��<��mB�ٯ�O�u�Z�Y��_�#�Ä�A'�O�bh~�ٝhٶ���4�2���:;/�^b	�k�455� H�w���)۬5�^�ٛ�����R��H#�0Pd���кA)
��j�8�=��g%_�}��Z|B�p?Qu�-����]/�[نk�2�6DV#�a�a�7�H��A��m�|Ck�c%��~gDX<o!���n]���5t�@�.����� �@'^�����ZE�Sb{�gBQ`���A���;VV)4��BՒ��.����C���V��g
|ߥ(�i��#�"Z]z��ģF����U���7pW}�'������6v�Nސ���k��;ϱ��#֦wt��#?;{��H��h'����93��G|��7J���:�)��%��G�Lc����̦,0߀�;.g;AFl�`n����tq���)@B��z?a�Y餪*���*�Lee���;�� F.�	�������)��xa�dF�� �����W��ϓ�dv�ӳ�:��J<4;���Ѡ{����~�Y�T��k�TvGx��̃)�m#�FZW<�v�6��M��UiX7_���
��o�̶�I<��S[�P����#�{3�/�j�?1��y��	w�;
����]i�j����`��>wT��<���!-Y��ViUծ�"��C��H������c���Qb����Ȼ798�>I,N���T�bb���=��¦�Qt6�{
^<ƃ����i|_#rt�6&{
r�0�Zv�����8�����Np7�K����f�W�x9��1x�ٵ��=t@��H$F�����얯f,���p�Ȅ�������A���_�j�B��������������T|u'dnz/�1�t��;W�@�ā(��>��5h�TRQ�S-��Cퟃ��F�g
�n�)K`ho,.uj���K}�J��klb%mi��3�����OU��vr�{54����0J���N��{��{�l2؀ŀ�z���cV��T���RῬ *X4���=�f>���	~c���'  �cx8A8t�sě�9Rՙ�vvn��Ka��!�4nI/!�7X�l�Ay��?QU�{��`i��ܾ((r��/	����F}8X�m��7��Hv���R�n�Vn9�_�=,!fff`V`���qN$ ��3��Cu��k�Z����Ͷ]t�k���7n\�۹l��ʈeH���K#5rM�������J���1��~'��y�tOUo������ݫ���}B(a�)��*_l �\30<L�5�E��"��Cgr$�k����,��@I2Q�t��w/���&]}p���L0�1kׯ�j�]Q��0�1��R��ri@,s�I�F�[�(!S��Bl��L^����~jgMU�����/���<��e��d]Ngk�<RnY|y��%Dͳ�:a�ѻ�4�ݙ�=L�R����b���F�|�t�;�	���+�*��%f9Y�t�1t��bKH����rK����R\R"���R.exA��<��;��p�ҕ��ݍ9��+��((ˆ9A ��Ii��G��]�1�)�&����!�Q��!�ݞ4Q�O0��ZQܶy�,՛�ȅ+1�tq���h��y�=D"z�i��$��@�K��uW�r�F��"BZ�2�';QgH��	���b#��e�ۣ��f7�~G�f�~]�Z���FJI��w����CVмv���������.0\�A�B.�1�����B.Donn���w@ؔ3~|`�Cb��PWn�����G�W'[?%�\L/J�z_Vwŏc�lx��0_u6��oek_����/�1��χ��D�H]��5DB�
��t�Y	N��0 �o� &�oD3a��(�}��M�|�''gyQy�`o���«��IE���z+�^TD(�)��������CՂ`�i'P|7�9�n/�_��m��r�]�]d7JEF�$i�3_t�v����p��{Go/��� ��W~4�u9I�g� �x�̨M��9Ҫ�}���g1B�w�"/`Ȁ�Ҷ�ЈĻ|�Kp-\�*�	�,_�V�ǳk��3��.ҦЩ��J�?K=��I��w����M?Q<+�}��������U��9�a����,��}E0Ϻ�#�j����u�zZ���Y`��Ք��;��-��j������eޙ�=	E=\~�����Ȼ@vp����B�_Z[[�_=���BTA��j�� ��a�N*Z���[�=� ,�c�2Q=�*���!���h���(&&&hT`UChw�atuu����+�_/r�%�,3Um��~��\6�ې����A8K=q��������x��G3��u�P ��.��= φY�dos�K�ǀ>�$�
�7�uS.��c�)QH�e�R�sɌ�����/)q �?�~WзS��b��ۘ�����x�4@�5?�&�������L�ͥ���� !�
�P�wi<q�^�7�hKo�AM3�͛7� �Ǹ�?��J���B
�������G�%�.�-��	�	�C����z|���:E��������Kd�/ӳ�� �PNNn�W������|��z 6����O��,&6��q��]���3�������
�39d�v�I�o1N�ۋ�}��*����`�FH�Ŷ}�Z�/������J_gd3avǷH��x����|��k���G5�F �b��htJJ
X"[/��-�a�'�w���Y󖥞���̛Y��:/���8��m��u�6 ��e锘����ϗ��7d�����}EH����O+�BAY��:#k��<�_�ēu�XnC��5�w���5\4-��/����z[2�T�77�J¤ȷ(e�l?F�����ȱ�G`Ls�  H�^�c�*#���i]���+�-/������}�>�[4�����ǻ���P�c�.͉����ted�W��D�ڈ���ӮzG�U ��8\��x�������CrW,`c^/wN(%��Np!��^���5�k�������@�[����Wߕ�O���V�@t�JY�7=T�pD������=��Q�	O�Ro	��c�2h.$g&o�ۊ�c�g�w0%�?��'���oD�b��e{�.2�n=�Xy�r4����P��_��H8L�='���׉t������,�d[<��$�}�����{�(h�|5����p����~Q<V�ݭ�~�k��n�c���2ZrZM��;���5ܟ���;7��v�����c4��/��Փ��W�a`���[�mv�X/��b;�e�A�Ò[4YHUt�M�����2�Q�{��_��*
�{�F��%V�ڞ�<��gg�G�B�V���"�k,�Ebܵ���al�\�qo_-�]��*�T��ޠ�'c��--�A{B��-�m�Aqb��{Lc�	��W%G�[�+�gY:S�a6z�>�vLF�X�3V�H�OsO;��#�f!N�T2�Nd���IΪ��CX�p�{v�q;�{d,�k�-Y��>(Vl~vU�/9IRZ�����m��l���w<c�(��#rZ6 ��^��D
+�O����(��
��<v��\P}��M�CHЈ�΂,�_kf�����
�������&6�f�"F6%��&Q��#XM	тiu���d����:���OD�ˑ�$a��������1���E�n_ ;�y`m���DW�i�͛ڔ�U��X�c��<C��>x$�3k�;g�����8���P�
�^�1˵I�Mn���pλ�������"Mޫ�zi{�� `�z�[��j��0�`ʝ�H	!�t��E�"ۿF��<V3�t��� g�����;d]ܜ�2�?��2n��2[sӪ�v�����lfn&�՘O�����IԲ�>��R�[ak��.��su�W(4p*�m��CH���G�*�).�/u��BE,�"!K1>o��gfV���\�Φopn�`��ux$���/����x���f�Qdy��ۏ�ܷ�s��@�2����f]�$�gl���t(>��`*n��r��!~8W�������s�T_jv#/[�@�isn�1>��8�*�����?@�PgR���]�Ӽ���rg�8/�1wy��u����̬g/��t&A��D2'���+���?�x���b�F��p�-�i�/�Z�fK��#�Mدlz{A�����;����k{r�,4�U��^�i��?O��G�����"�k+�(ޚ��:�m�9�:��W�uH>���,����݉��Y�J+�a/�*C���k�6�v��n���������]��^�%rY/�����Z�L��3�5��<�x$���8��z�9�ʼW�e��3 J�ڛ�V՘����3<�\(�5���,�6�H[	��\q^y�pY*����$@p)jml!�JTQ|~��ަy��<67m�W��iN��.��JY�@x�����-�?�����OᨡQ����0=�@p2����w1��7R�������8����-v�7��ʅ8�O�Ȧu�=���a���A*�ס�MG�E �L�m��V��,��j���ƒ/s����T-��͏��x�y�j)���2���^����%+|�W����@�v�B��6!3�!�U���,Fi��)���7u�٤]ʻ� r%"�����Nd=�0���J��kZZ���&v+k|�+7,\���RD����љ��0�m)�b$?V��������L=]i�7�j�X=w?o7F$��x�U�eTbǕiKE��Ґc-Fzk��+�N��uR�������5��p�m�72'�r$�W�XOʦ�Z�����+0�N�&��ۡܝ�)�R�f�w��3{FZ�����֕ɼ*A�"?���i	�m%��ȑ����0y��Yq�9ލX����͆Ô
|��s&��:��]˭""��c�m����F��H��z��Bぃ�����R�
�ي��.?�V�[���F�)y��*�����
�՘\�pݪ��-��dXYm�dO\�bUŷ���W4s���"1CW�#���a����Q�O,��\+(�x�""����󐅰���&3f�_�)D,L�[a?���PU1�����C�rzH}!������Q�
��o؂	 ��e�oH�0}�5{���S�]b��:PD}8�y��Y�qL�Klo��I.��j\�t�ȯ7�G��1)*�~d`;�5!��'���T�d&�U{Dኼ�7{¼G�!�ԫ�����w��N��o���u��\D�d��R�⣎�|���jq�+Ĵ̓��s���t�RN%r>��:3��a��o=u;X�%�·HYb��j����[V]��|b�؅��C���5EӴ�*Kc6�zg0����~�p�G�2��*�j~9�²ﵘ�)�,���b)υ�<����S���m
��I�ǶJ["�J��~����Jy���f��fӌO���)�zHeZ�wUߟ��E�#^I�:���c������0��O�O�gu�,q�`J���X�	:�7l���7���"�GߜR|��<�����o~����ŀ�Q\`�8��A�0�`:̞Еvݙ)g"�޺��0j���W����f�g���/��(J���\�@=�e�K��Jo�0u���R�[��w �yn���E��W�<��󄄨��V6P2�������Dk������,�S�?���f�H+ڑ%P�SM�j���j�q?|P��U�:�O�(8�˫#�8�6�/켌�\=> 	$ڇ��.�G����)HJJR�s�j_lQR�98�#�M���\�22�� ���<��UUO	���gQ�I!�}h���{!]���@�Ö�R���0}�K�������+W��m�� �&+���+A��s�;c�����id|�\uļ�E|x���I��-�z��\e���E�_�05�����ݛ��rAim̄�����C(;������+�G+�xv��u$�8�,�N��-X)��x�W��x	oo�w�����@nL�&z¥���uj/��_�7@xי���s�H��l�%��� ]���S�v��>�����Z���EAB{����:�5��v�ih���
x�~�J�i:����%~��x�Y�	&��	�~^��2!��5�_7���Bj��ȓ��]�'{D����y;�. �rGnhُfln�[���5X7���kI��N�]*�V I�p[e����Q��A����/>�߽Z���=��
��Q=M;�?�����qQ5M۠"(�J%�H�9����3���d$�#�P2�$I"9�$�"90�9��9��~O���w��ﷻ���8�tw]UuUwu5�;q�[|6�)[�7�!���ha2�V��1_k�w/1�Έ�)f��))п���c٧�@B9z�;�c�D-�g97~+�wo�i����ЍAo�Wp{%a^c.��r�GV�
'�L�17[�N�^�0�~��EO�6��^Ͻ�x�=.�C: 8ͭ;y�L�{�쨒by��DSya�B�$T����*�h�10o�(:��`�K����h�P�)�7�W��p_�;�z8^�>�$���}:Xp����X�XpQ�ߴ���H~��Rnt���:Y��8�g��5T
n�AV"s0IV<�ӳŲ����������9t��o?�!��F�$�~�FU2��'���k�0<�E'E\�=u��.#��\��];ꄄ�f�=��x�B|P�dGY���fY[[�HOO����z�iڥ���j��His(���I^EFq|�HY�3��ɋ��ee��ͫ�fp��gΤVV�$��[��X����  �K�W�{��vW�:��Ν?/���+��T�����6i�]�P���.�ф K��`xx�$�2���tj�HZnɏE�x(���e$�]�x�ů]�$E|���.��˗/�WS,�~x�d��(�1�*��]s�'���R�p�m;�#�M��"� `��+%%�{�b́;)n0N�++�h4����ϖ�N��`v��%�0�N>�]��44���}�+�b���cڎph�L`�K�u�n ��/ǃH!�XxEE/����ND�0":;;}y��3�lf����w�;��������EW���gl�>�L�����}K@�*/��§�����!899����yzzJ3�t��� }@l�K,!���À�H�
���dd�0� �R�An��[Ź��
P}�9*��p3y!/�X$3zN2(��L �_Xh=S���5`�oĭ˿���
7��P�O]Ӂ=�Um=�)��M��.� J����`�߄)��ڵ�M+�C�@�����7��u=���ؘ�����^ZY�L
H��QbWJ.(ࣦ�f7Wb�>%4��Us��2?x���s�1���U���
���j�������ɵ��6��W7/>���[��f�-D`C+VV8��L- ��顱��Z5��y�F���[��k!���/������T�_�����KH����x{{�]楣�{]t�:/
�J��'�OΥ��K�� �}�����Z ݇��q��+߽�
����~Ր^J)É�Z��i?��G�����^Ⱥcjj�5�Q�G�V���=vopÓ��6�22�tw�]d.���m�׊���Ԍw���+Y�6����6S*
��Ћ@�{h�|���6eY�E��p��=�t�j���E��yJ<�*i����B�3m�W�������H�����=Je���|���3����E����n:�ڈCy�+�L�Y^SSSJa��.~�}V��� e{�6CYɹH�y>;;�UO3N�@�|Kn%�W�kz/��$`� ���Y��ӊ���������9���&�����w&DgSE=j����OM{����~��.j�s��Y�Ą����<�dж�����rGR��B�Z����`ֻ�]��֖^��;FeE7G�dޭ"����*X�jCs��Vb�}���(��G�ᗑk)�#a�D�K�Ї����]Dˢ��mO��!�2h�_�����~�عv䂂BCC}]���6|�Iy}౱��66-���
f�7���P���&�~	'(i�uH��.0l��u��r��]y���
��f��}zVPXp�̧��<���V�4<պ
�Vj%�)��v�aQC�V=��ߝR��O��s@l/SG�u��u�J���'y���/��\�/f�e�7��7�k�t6������[!AzԀДQ�`�gf]Z��n��_��9����n��������EÁ��N�^�"�B�`��u���'�����؃��E����> ������)�������������� ��'���j�b2nTw0vM{�[b��N/�4����ù���:ӑ��\g�L�Mfx�%6{<7��$�q"��F|��*�J����%��~���P��� �x����a��Dn�&�9�Lː-���OeM�${����T�Y!B&	�EV�\Il.�v����N���ľ��z^h�Þ��97�]��D��UW0Kr0ʐ������~���j���Z�{ \���(@1OAA�:	�\!!!�4��"nO���b�����dve�
0�<�q�!40�<l�L���u��2<�� �j���
�v�	G���h�N��O�Ү��Bz�_�G����W|詝��p�t�S�NCp*�q������ۅcaa�[�t�yWj811���[�r#�D]!��8�g������
٭%)^T	����"z��v�Q-���\yD"H <�U%9��5����ߟ��6N90�:����/�+���;��Pv�ݬx&Q�r��X�｢�6#4x�*�'zFF�d*+*n��)ڱ�47��^��@��"�ǯl��ͷ��Ѭ�Dj����������͞N�Zj)��3iĻ�1�h������(���5]���#=g�1e�ؖ��$Uϋ�*1c5�k=d^�p��oD$�X-y����̯�7?���BW�[���c��' ���焊K�yc��D	�7��W�]i.�E���:���Yq��a��C97���2V�Vȷ3�b=<�����v�4����x�~�]�|���#( z�Z6QF8U�\]��!�]b�)��m�++��"5�b75㨑i�2,i ���{[�B`PNlmk;Lq��H�y�ϼC�;{�(Ƭ~ǆT����q�A�����	uc(����e�:��W4���[2r�۰��R^�����4���
��^��j�ܵՖ$�/��]�2�
�s�M����Ö}���u�W��$:YG6����Ea�(G�ޣ[w6W�m�}9kܶ��Za�������x�G��_f\���K���7Rw����/�R� pV~�H�_� D�̍�j
NEES���i�a�|Ģ�c�;8~�5�iV9���R�l�ֆ���8OsL囮�Sn�h	��G�F����.P_�{�T��v���~=˫dn�+}?f���K����e~� �ݮ����d�wt5��ۆQuQ�P�g-�]�qon����c����
ij�=D{�o���w<��^Y'R��Q�=�3�gBF��bz�I����ʕ�B�Mד��,���}�VX৬��j.��r��!�:��'d#`_��@��ȕ�u�>yD�q������.mc:a��ǒ���VaA�P}��n���W����ss� ���$����ȚnkZBƨ������S������sG#6��@�/�&��n�p&)�2�*{iA��X��GJJ
}�
�=8���#���
����B��3<\�qѲ��]��}zA�3�AYU��`%��|YҢp�&���E����I0� �$ݣ�"���mO#��b��jRXFE�A�ݜcŰZ1u�c�W�^�.����T���w�*���0������nV��˲f&�6(a�"8�����f�r۴�J!�	��=�УlyS1�tA����="�mh�M'>�W�Qo�ӿ��'�~����{��}������`�I��Կ��F
�ኟ�@�V�$�8�,M����,�����,��L�ڐ�"�X꿙�3�gl��%Ľy,:���ꯆ�!!�ݡ��� "bΏ˼������j��IX�^�`w���)���H=��	�	��E�^�n#��+���h+t�OY�,�_K�Oury6y��Lt3�B>DV�[�8V0Sg�[b?�w��X�.H���R�W�%A)-�H:����~K@D <v�}�C����ksW`����0�S$:3�9�B[����ٮ�D�{*����}P-�,��Q��ʯ��D��0�mع�+�9Ϗg��H�fc��lmI:`(̰�[U�c�����i�"�Gg�غ��mAR#;gf�-��H��� ?�L���
����u�E}�@/٩�S��R�e�}��Q�M�,��3k�R|���O ���lݹ�{̧�����ox:>��o���iWJ���	w����yq����p>aa�Y7ps)}d'�x0��e��Ql��ˀ��|��2��q��uC��^����O4V��b�@�>��3��@̼�@?$��������X	0?b_;[G��x��=��i���(n���{;>����T~6�`ફ��QFw��r�-����d�{�a�cQ���rི@<�@�Xx�,bZ�55�,1x�&�����qh6#9��z1� xβ#V赤'��A�׻�qP��XO��ŕ��@PhYޢ{�u��P�T�&�!$�3����?�IOD�~Ry��Wh���Q��,�F�yhN{�������f�e&P�q�9_3KK�7��ܘߥb�byY��;:::\cG�B�o��P�j��g��0ν1��9��W��%���m��QO�F�]<��,^l�e��p�3����;���)��nqwa��[\\��4�Gy kW��(�)���u�N{uY��8�yv�pKHF��PoY );������ĈFĴ�ZEyy��;�<wd�B 4Y}�ށRʈ��Vo�;��[�i��#y@(.��gt)0�h�wV]V��@?��o��_vF�@�{���m��Π��7o��\(4Y�V��"���x���Y���aj����C)G��?�3�<�-7F��
�q���T�j}<F0u6ǰ���g���؍D����%@��]�̀� h�yg�7B0'B�T�m�"ȟP16& �������`��%ß�����QDu���KGVUx=�LUN�9L�F����v��Q�75���܇��G�~A��L]����A^8��3�V�`���!�������[�����Z%����^���Du�ݳ@ ӌnf`�F°ᑯ�2R�Ү1`�/�8��՟��#*G���:�)|���ZeC� ��=�����ɛ�"�,_�h�E�T.t$��Z���{ݺ$�����x�Dn���f3ݗ�/p�`�b�R&���b!�s+�"�}�y�c,���	
��W��3t������qȗ,I�'^ 1#��@��EL{�� �HT�g"�``�	;���@�6�����Z��BV����`�a	�ec�k�4�#V D���w�ǼP��YJTz���L?�T8�d�(?^�ě�j���qi�����H�9A[Bo&6� ���%9�c�T��r��x4����=�"������?1���Љ	�n�_��L�'�r`��u/%�H��$n���].��B$Y��F=�|70tN��"�W`ޅ�A>��;��X�y����[��	����KNe_�L���Rz�U�7��lB��d 3������X ��xW�gX&^�e|���guk�]�y^��{)�©ǥ��X�o�f��o̯��ɧ{����|LWL�J.-)q���y�{�@唋��@� ��3�A�jia��=Z�����aEww�Ej��_��|���Li�ۦ�P(d)���M �ں�u��r��[v�/Z������^f4y����Ho4��K樘�
�w�n2��n�M�+L��bRrK�RU˓�F�� M<�:�sG�?gmu��r|�2�Q	��o�0Ǟ�+bt��\�ỶJ��]k�ύ�5<�F-�D�M��E��+���1+q��;3ƇE��� {8�{���a���~��Zz� ���~��ӿ7�8�~�F:�1��]ч9bhu���x_�ǜcV��ǆ+|R�}3P�%?77���$vy�T��jտ�7*w���j��U�3�<�����\i�!�)tjd�+�)�=��4+�G�	<��d�f�̢)����f��U��X̪���1{d�g�m�}��dI�n��鳁�]d2���{�>���1�z~x��QE���n��]�O�4����g�7��Fy�k\������v�ü��Ύ755ٍc�J���&�ϓ�^烠S_�,��C��SFRw�����L���uCz�J��˧Ó��=1�����;����^p�9Ǩ�?j�'�{���[�zìC
��]�*	�o	AW����܊�|�����\;���ӱ�$ױ\r�@�n����.�n�N!V?ޯw��M���@/Y������vq�|���r�o��)Z��h���U�+��Q�y�+�mQ�+N>#���++�AC��B��n���d#�ܫ^DwYwF=��j�Z�����؞
�������������y��qUL3���o�?����sȾ�i�cƥ{d���^���Sl��n���s
vV˂w�����Ƚ�oyBg��u~���fT$��ؗ�(~m��xj���L��<G�v0U_��ͩB3?��(?�ۙ�B�"�͛7{{{�zJ�a&���i��%��ٳ+Vl�W�0�=jt0��TVnS�ٙz�4�F�¸$�gʜr<�~�1��L���.sN}ɲ�'�������a�n�a��]�S��0�J��ג;���Q���n��-��]����ݩf����μ�85Mj^7�[�WiL"�##>�߿� ��� W<=9￞?:
���N��B$�M��V��A"�[����t���O�+}�h�������w3r���P��}�����+k�q|��fgga��vo]��6!�\��宋�&�i6H��Te����c��o%�Ku�>�H8g�شvc񵢕�xQ&FQ�ݝʘ�y	��,�uM�����wFJ~�H>��m�MPH(rC���0K���/Ow0Os���L�kũ{B�����8;t�Vɵ;of�I
m0�U,k��%_��L��0�so��8	�t��>e������/��V'�p�d��-�����=�L-8xC�ESs��G0�u>�yeӽ����<"�[�����?]��H�k�9�>V�.�����)�����0B��˗��\���<x�}�/t�F���
�G"1I���ͅxIE��k9��>�Q{��@�.����s+lg��@�I�3�gɩ���/d�u�b��>���/&���q&3\�9�8o;\X�k�E�А����Z5����h�;NN�?���o�uw$b,��EP�����7a�Ű��ߏ,]�m�M��C]�]���j3$x�u��$���`J��A4W1�΁�H���ە�Ͼ뙷���E���4455�*;,�;;;yTȽ�}��|׹l���yU|����0�B�`*ƴ]9M!_Z�S��_�f�LHO����+���Ƅ��V���+�y��h��s�1߆�C�n�'''	]ʍlk�Ɂ�L9�Op>?_�+��UV9x��Y���)�.t��&�`�!�b���]�RTs�������	��8����c����ᕖ����gf�310�G�X6y~�����=����:���eG��JϜ/���J�8��sK�X�z��C�|���5?m�3��Nt��~��=�H�f�c>\�]���4�)�s��c��V1x-��� p��+,�=Ӵ�I�x�ϑ,���v�d��Kv����$��_o����{~�!���@~�Į�`5���L���A[*�'K �(��K��;8s.埉f��;ք
��}҇a6�K���x�&ċ�����Ψ �}_��W ���U*�y�`8�޼@r�)���J�q�y��_����.����7����l���i�f���e���3�b6֮S1�g���޿�2��_yS쵍K�o�q�u���#��{Is6�0�IArh��'+I��-�i�l	��54Pߞ�r��{���ݰ�����g�w/�|+���	�Eccc�M����L3x #�����؁ϑ��4=Fc�pI9�Xr���=!��e��{�~�̶}R�/�o?�߷������~�O�gS�8O�F��UO��=�_:�����������CTQW���僱]�Ī�4B�?hHYh���5'''A��~'������w�3~��Vi�g�z����b�i�]���ո��t"�;�PhHȌK�Z^Wbq�Ư�]���7QG�(�Ra
���W8Xg�ð���;�4�$�67���*�I�(�����H<���|�۷oo����&Y��L�i��5�=~U�B��/����bBT�Z�1*��u1YYl����AvVn�=R_�6�f�>��t~i)��K�}9�9��ȍ��T�G2��{�ĕ:���Y���Z=��U�d����#�p�EZ�v�G��i��m�.ķ1�!CBB:�vV��y�f�W�9��W�|�IP�$��^92ڂ}B9�v�?w���y��.��A3��t�G��.�#w��gm�����&�ĩ��J��%�hٌ|L:��}g7ջ��"0��9���[	x��y.#u�ܗ��)��\�3���:$e6[жW�?ǲp�~���0�={�C��0kX�Cs�)և�}`:|�uN&\�y�<A�R-|ܓ$�c�1������O"�-+2�+!�>'���9�9OkE"�ͣdIR%����� �SiuB���6�(D�3]Fܺ��^��R��a�j�%Ϸ��p�v���n�t�u���٥n��:��nk4��@������o}u��Zʹ#�-u#�g���f��Ƒ�l��;x/QOkb��� ��l��<5�gѓ�*թ�6��| ��� t���/4`�:�3��kt�٥Y�#xR��6_/�O�ʓ�Q�1G_}����ma�-�9��\�˨��*T5�������{�͍~��?5�z��"�;�춨?#_db�z'	���1u��	�!���Yv@�:�19Ɵ�D��-��֤\���H�҇"]h�
���4��O���(�`M�_�e| �S�^��(����0X�(�ڭ��d}��U�驘��'��T��8͡Ƶ�_H�3_ν�R�4s��V\�mAfA��^NO
���P�"Ab�_H�����5Ar�^6����k���]����¸nN��?�e�8��#������NC�� ׌����T!�R���}��K�d�˶c�� ��>�s�	��9I��9���.v䚜����_��)u�s�0��ԟ?���<Ir3�Q���^awg:"���	[9P�Q��Ŷ�6뫖�������� ��� !��a�8���
�|�T����uT��L�^��:��ź^�tfn���؆2F(x�w��KK���?����RkW�7t�z_�ӛhRg�Yl�G��$��J�h+�E����\p�*�y�|�Y�5n����uHT6�x�/��Gc�_��O�=����(`�2�~`I��V-hc[ڤ�ov�?d^�2=m��+P�H��:�n�׽p~_��^ ��ζc������N"�<�H>�~0k|b�h��c�zG���UÇO���D�C���1�X�������V��Ns7�v$�����ǥd�9�@c	���v>
����QMJ[#,**m�������:��v�R=6�Sm�n�9���Zz���D~��v�$�qt�#�����ڑ�P�U�1��M�����~�tL��G ��/��-��L��4��F买�i���j^9�����ԫ�s��&�J-�ЂR%D����6މ�R6B��c��?x�ݜR�����5�<�`]��gR�P���������޴>��B�����÷S抭�B䛳9NFH�5t�5��S�Q��pc&r��)7l|8:M*o7�seu'�t�}��_6�p�c�~G�\^R����f������ƒ*�prY;�2���"�#u�،�W4��%:^���d�(�ɱ��wdS�U�V '����<�Uf;�]�<�tS~�~���E�4K��o�p��f����&:PH��U� DJ���X���+��0���*z��E����7?[#o��%z�ymq]'ʮ��]���v�Q�9��	�-�W�tj���j)��DE:w.�5��K��������a�l=G��r�ށX���Q�`?79�9<l���wm8Q7j-v������퇋ٸ��?�d'hHM������E���7�b��N��10sy����G�X�M���*�iP�XV�l�.��Y)��j�mJq)qq�vWN⤑|_�.����7��>XID����.�7F2T�w&��ǋ�64�; �����Z�l��y�-�j�:Ue�+�V�Иa/�w@57G' i�}���N�(�j�*!L�[zU!��+/5���:
l4'�#ߴ��r�Lf��
 7p(cl�p��""4��*��<sD`�g-݈A�2vޖ[�8ࠍ��!�}y%Ɛ��"s��wV'@Q�5g�l�(x��ۂ?��¿

9��{�-��m@��s�P�Ҕ߭��j�5`u�R�z��[�l�׷��9#xpp[Y>��W��vϲ~��q�	z%w��'G��V�i��qД�ز�i��'75�q���r��7�Q�	e������+�Ȫ���<wtvK�įK�^q&�Q��z|A�2�Y]�Xl�?�F��$�B�W�Q?����`-��ￌ�d��Z~�/|ZWv���95,���M����|��`��vwy;����J�ƭ���}Z����s+/h��nҊ|Yy��������&�<݀��W����V��5��Y6�7'Qd0�x����uQ�K�r����X��ͺ2������HT�Tqpjnjn�&�1�
n@a��J���#�%�������ŷ1̀l�_G}�RH~[s9�C��,���l��jr�����O
Y(�1lOd�b�h?mݍ �;u`�U�-��{�Id�MD���Lv5n�`���1�Yy��%g}�Zܧ�|�}W7x��I���.&ҼC�R��M�w���^�>���[yt��ݑQsIbk�u(���Cp%
���fT�#���h$Ms�T�ݰ���:���~h�$v�;�~�~�`d��慝�`L�;U�3��|���Z�l���η%9].���U�'�lϜP}E)f��]ۧ �_�<Q�����>��1�&^$�!/�[uq���(	jJBח%/�Y�h?���r�C6�q,�>�We>�c�0�����ӥT�ܾ~}r����s�U�卉E����
G?�UD[�r�a]%Μ�����U����Q�6��b���Zb݃� ����1���c ����&�yN�_�n�]P��7?���nI�5�]�˲%�9/�߰���T�ϳu����x�J�gS���9@�eCΪ��r���wYܯ�"M X,ԸG�h��3;X� X"X�$����[���|���un�`��}I������a�P�oϚI~)$>S+d�nq�7 �������mh��6���,P��uam���y]c!�.�>�E!"�ɭT$�Ϊ��0`�Q�Y��0�<K�u�X�Z!�mAʢ&&H&2䵨\q2�7q*Hb�M����&�yw7�0��L,��7���evz���{(CT�3��)d���*˓@U\��~X���b	����D3��$ !�x�wv�Et��=F��Qt�Y@ Ae�qO�c��_(P�v��F�{m`�ԏr�^H�qw7������i�����B����x�=P�ʏe;�r2e�A#��RH��q)t���li?���дE$��[ZM��QɞW��g�h�·Zʃ��}pP�w5�:��48Y�lZ��h|՛ cع�.�����)i���a�M��'WQFqްm�J�Y'G{��X��y���4M�	Gh�_(�'İ�Ъ�|��o����Ν^Tz�:0��5���;0J�jlΚ��;�������!�w�O3�g�����ht1���b������$UR�>�7:1h��3�m�9���Fu�f\H�Y�{�RM�$=��;�,/5~����)^U��|��3��R�+�~��(t4n�/��d*_:��7����΍�� �LŊB�a' �tz!G�Qnh�����f����ȫ�c��#z.�.��|=F�(0jU�3JC���Ű.	��k=�����������W�5N��g��.<V_��u)�i}�k�'֤����Ǆ��po[�2Yh  "@��K�퍯CC�?���=$#�z-;��A9"H/Euj��L�BcY��;�.�9�E��9��Ft�A+F�Y1)�@E��d��_�&�,�����x`��e<b�����S¼�œ��ۏemp=V��FJ�0�\��m�}�lM]��U�#�f��F#/����b��fOޣ=zM8R��3�>(�{�V���GX�
�������T?���C�4�&����p�c�P|I��@���5�����'\�9�u��H���עQ�̸��M�T�i��S���|�x��tM��Λt�n����v3�esV�@8/�)�h�5S�d���M˄`��>��y:��PI����]ךz��/~����vm.H�ߛ7�.�u'���1G<R'�)�AE��W�$��U�-����)�B&�X|Di!Oa��H�I�JE	hKԛU��h���Z�kNRe��`��Z�$W�zq����\���m�'���ؖ2��S��[A���&*�ӑ.B��9���H. PW�߿4�QJ
�F�3;x��˼���eU�@������U{ɀX��X����ɛ���u���$Ͷ[�V~��7XQ*T��l�T� �Z'<�#�2��.5b�'�;|�N�ȼ3Y���j
�f��X�r~�@��3���2��d4M��:�����=��~���?�?FE��BJ'��'g�<ēuq��jt��!<�c6H����T����'u�FP�}H���q�
P�SN�
>sC	�{M�c ْ�e��T_Y-':������&�۶%-G��'��O���m6��fX��;{8�zs�����G;h����=44�|�o��<ړg\i��6���9Q`��T�2��|/_���,��q�5�krӽDԐUҲ�sD *LF:]=��%��0��PP��w��:'>X��aۧi�}4�/��S'q� ��9��*��.%�&�\���.߂�Ǯ�b�!���S���6��g���P��hI.z�ˮ������9���L+��5�f*m���xIu����?f��3���}_2��L�3�2jH�KJJ��Rjv� wo�\���^�}*����fҞV{�X�H[�5����F��@id���F�{� �I��T'"�]ʽv&�[�U�;=�n�DhdC}�h�$���ۡD����Q�4o]��4�M㻴���+{�0���K�];Uf�d,WL�`T�R�З-����n�іLװi�	�	�����^yi�UV�$�sE6Y��M���H�'������@�{���s`L�c��Ts0>	�6�Ph
b52�A�����=��H�1n�ݥ�����m"����u��q߻�J?K~��/+����-�VK;zO�V{z��P9nE�h��(��֏�G�s�CHq	���	!f(�2 �o��V.T�Dg��iYi�%NH�<�٨��Qew�7c�d�l��fj[%��4��;]�C0�۩����K����r��jߠ�Q�¹�����4���f�$��%KB��^��Ɋnp��T�Ǡ�����}���W+ 䉾��Q��1��K<�6�=K� �7hA���K��}����˅S+V���+%��G���7\� ����J��I�/�����[��:@h�p�h�U����j�L�J3N�� �$N��=�}?���̖)O ��߁�z3�%��gj�~��l.d\�f��ү_�����P4�h�ڝ:^R��z����U���(��0m{�` "���M�3��`�.�b�P���zm��K��W�j,��e1Q�G�+�A�]?{��m�ڃ�k��u-��ۜ*��)&-p���೐����$�ܰ�,�j�C}#25�V88pM
K���ٸ�?�#;V�hU:~6ǴV:�k*p�\S3p|8���e �W��8{[� �$_��}͓}��E psp!ʾ�t�Ͳ<��R>����z���o��w�Q�-������U�Ş"����#��ܴ-���kz�@��&>�8�	$�֎y9��ok������h�� _W��+*)����)/����[����J��Tȵ���-�����k>>����%~�ZA3u��.H���u�~������[���㉭��ռ�u�q�����Jaz��I����6���L1k.��6�^-���(�?b2�ߝ99����<���E�c��9�?2�5$���x������/� ��z��iT��О$#3�rU:cy�%�N{�>Ѡ���j����z�.3��m�B�\%�*��m�bqMS���)r �L��!�4�YX Y�I���`IO���sK�f�@��۔_Y���ާttt�S�;��`t����1����N���o	�+��ST\��%�.�yr���m�ۃ�ɳKx,}����,q0�1��=XC�:��fk�C1c ��׭�����z�Ay��������\�D��6��A��v4Ĵ��ڶ�+I��q!
~�+�X������ڙ,Y?�B�Do8��-���`�
�P�YD�@�,d�W̪���c6 /6.�b��ӂ{����BW3���ϻ)�V�[�� �\r�42�<��:=)tx��2@U�ƞ�B�Db�� ��	a-�p7����k@RX�Wc��6�v�i��s���ɫ�B8����̘���-��lj8�!�Sq܅��!���H�pi��A����a��\�C4�����Ų�X���!����I~���O"Gǃ �<�{�钾��n�Qr0������~[��up�S՝I�H�p���ng���Ǭ1P�@¢���d�h|ۂr9��7�� :`_d����YC�9W�hS�S����R�	r#���ec�tftG�J{�������w�A��F��0YVU$���0�R�뱵+r�?<$��¢�i��=%��i#�[B(�Chh�Y� ѽ&	�s�`2"�B&�+z'�� ;�&`�m[���K
�+-6(�r� ~+(��
:�*1��@#�U�ǲ|�N�����p�� �����J+a��E��9oe��
M~�z��'#q��/i"E���Zc&�i�if8?�C3�� ��?�F{<5֟oM��;ަ�|�GA=L��������z��Lk��$��Sph�Dr@S9�gC�E1*��n;K�Gh������Z,��Q� 3�Y�������>.�?	)rv�)MKw{���BZ*�6����ii�J��VJF�	��[#[|vԵCʹ�&Zko�7Qo���z��ik����%R��M~���Z�u�ߦ���(�n_NțƱx¶K/����M#���&	<�E�����9�J��+�7���&Jj���Z ���n���nB���1�q��qu����rW+$�n���i:"N��d�ZA~�K�-�0��J0M=�63E�4ޕV�xa�b~��õȴ�
d�� �FZ������Y��ЌnK���^/J���S��Ē�\���v����&U��^�\?qП6f��PT����_L���,$�p\�D/���q������Y�^�鿈��\�t��S����9BG���]:�b�M"ty�?��B�J�v�mi�
��.R3W=�}��rN��5����^Y*�j���h
@67��)�~�q=�%"%(�������0���2S���w�iL!z�#�+w�������R�����}�Y��j�f_6����Xg��j z�F�������?!~P9��/t(�_����;PI��o�q�K���(Wsk*-�ݢ���]����R���@�FB��>r�>�z@'�cp�HKGB���d<��l��i�J.)$�f��%	vP�?���A��5Z�xMO^���4��N�LWY�__g�l����qZ�'��W/'#n�NS��k���K��d_�ybNz�?t��EWVC��p ¼�?���?���?���?����g@���N큚�D�bm�H i���l1�����>�P��m%%�}�
�~ n���t�Պog�FH��9���Zq�u�Y�L��L����z�6)1��	���iRX����1��J�z���E�����~�\�ľ�dF��Q��K�jvKɉ�]��j��~�Xt����=����h�Ց���:F/f�-+�ܾ�k�me��h.�%&&x�-�BS:E#�j���do�)������M3�?�f��~�	�"&1a9�`���su!�n8�Ӄ�@��@��@��@��@��@��@��@��@��@��@��@��@��@���CA)k�C�2�`��S�q;�g�!�?���m����:Pb*wG
�;��H���-Mc���mZ5����e�^O�ݗ��8����]Y��P��5��֛-��	���;}�(2�sϓ��Aə���6��2m^�Hb��]�Bқ��o�J�t����A&!!!�;��Qi�ȓG��^�'e��\�#���X<��|��o���^ �l�2��ԅ��SP��=R���#2�ۺ��6	�&nyv�md��t��9l�e���&�r�����<�r�[p��Nv��a�_��FV�-w� ���C(��p��|ˣ��+��_�ݴ���������S����$�]�����3�v�n�@(K�_�p��Y�լ[4�Rw@���>T�}/Kr�u��k�j�[�����U���,�,H�5i�1t}9B�z,Tj5��WXg}�|sJP�sS#����>bA�4<8g�Yg���:�K��g+D"_����aǎc�q�q�֖����\F�P���S�
��9�e�ڪ����m��9��'�H�Bw�dV
^ ����s�l܇�+�P�R�ݤl���ѹ+�Ji.m'bL���YE����p��b�l�h�]&�o�W�!���'#���VRÇ[�mU,�Sz}*��ï�i�J�k�{p�Μ.�m�����ݢ$��Na"�́O��?N�3i��d�q�׌,{\�(p6tht�eBBBu�(z�q�\�pG�\^�9q��	ua�	G�Ոj�s��Z(��}�u��B���n��fkn�׿� l�����o���~���h�z�FTzw"�;Sd|}<@�OF��qx������p���_�|%����@�w��ǸJ�G
���rf�?[ 
Ed��t�WD4��U���yɻ8c�"�����m��UY[�i�DB���K=��5�?�l��o$}��G��q�ޫoq�Z8n�z���fr8���vkw�����۫j\���guj)��R�C�F��&�!�4�
Ѣ���_����5rjྫ*ؔ/���)�M��H4�gO�~X��Y!.,�:����c��4�$_[[���Ms�6��=T�	�n�y�Ǖ�����8�t��s�l��×�^r;Ǔ ��� �O=P5˨%��oE�.����4��25���/8;���|&Z梵CV�ߵ ��|��U�}����mB�F��>������m�zl��6Ҡ
�e�m3p�V���א�-�x���ZG���]-��Ȝ�Z	�R�(Ԅ*K���`q�T���sͻX��z!Ii׍/��,�^�ʹ�Mo)�ާK��]�A�[>9/�:n����T�J��J1J2���F.V~�2����`ۣ������$U2S�����i��Q�S�����x��*�^j-t��t���	�{������`�Ō��[�}���������l�KK��� |TP1�����L�j�햋E���7��OU�͸-��N~����'�6T��B쑭E�b�~Փ\4(��h7��ܟP%���`�_���y &�����Y]g�ɹu�6r��cL�I���)�=�����u�9�.�9.j�����c�fi�C�y�BB�Z��}P]Æ	�"�/��7�/���-n�� x
ru�z)��O��o�$�S�R,�#NXZ��B�9��6�����b{_GEYC�pF!"ۧ�IW��p�s�r)�&�L�s�3nE)\�6�m��@�s��!�O��c�.«WK*�p�I97:�=s��~�'����<��+�z�_�_c�f1e�>�n�S��uf�GG9��\�W�@4�fQ��F<`����e-En�WK�/��L��>T{���ث����������#� H��A�R�+��TCo	��"]�w�J��I�5@��B-���N�;3��3W�y/���s�^{������Y��F[Nz��D��|�b69C���G%�zz]�cu��R򓍼�x�k�~���h��`�yѦ٦qp}���^�j{�q���������缧dՑq���w�?�P��T���\�9� l���|5f�̡���7� 1���(�ԟ�����[Gmw��j.������@dZ�MѼ 1�����0JA�����j��T3c֐a�Y`g�g�o\�����Yz�5,�Y#ACu���E	E������QS��]��h|�s�Ƿ��TtX��]��X�՞(�?��z�L&�`G����o{��>�g��D� f$�>��s� 8�ܰ �S=A�J$���6x��q[2�U�1�Ñ��ٸff�V�XY�bW:�M�d42��͉�8��=ؿq����}mm���Qw�Ӌ����;�o��P��董o��?Zb�6^��M7��J<�.��d0m0���d,�}R��Ҙ�g�Ѽ��\X�(�횢�#.�G�uaC%���rc"ڼ�0~�t;:��'����\�^Ɨ	�؄���̉���f���H�U��Ő(��w�N�;��V${�y��c��ۓ�����tJ���8��No�_}c���r��|o�E�����eiQn���k�@L{x4�֭))t�?���u�j8���S9G��@xH��5rz��[���#|n���� &�s�M�o���;��:P���~��Z�O�4J�#��8��9� sl�YA��wNRE����kd�G�R\��U���b�a�>(]���upyvt.wH�s��)��"@��fNSΗ�)��O"���o yc�o�yjg� ��,����l��b�D�O�S|d�<�&�W:E`�~?�v�J���1��d]%�^�4;�ͻ��Uꏇ@dF�5S�>���ט�=$��\�i��)�D�L�	�By�¾�� ؃m��S4�-r �C���ClOR*�s���=C)���]jϘ(�<�����r���\Qq�Xx�n\�������G�����4Q���t�T7Z����b��&��֖sq{$9�	�����A�!��hرɜ$A]�{�2g0���5���0*CR��7����Ӗ�tzڨI�5۸~��q��T���9r�&���d~�������7�~@^���Ɖa7z��Yh�Q��j8�A�P��*x���EB�`���;�Z؏�Z�)ۄ��s�s�(OK�˟��D֣��_�gى5f����sF��Q�Y�����g^d�:|����:�>^��R����½[l����&\��3�h��SV߉P���IK��7R�)}s-}5>e�Qfڑ��X�`���X�$�V]m���V��C��o��.�%�fa�_�|�����gO1�'�H:y�K���ݢ8��;�ʦ�2T���b��q�)��'��Q��͜ɍ?_?�sY^�>�&���{W�9�.�vQU�V�Ʃ���%��w6&�����e#@��7�e���^8'�ᯢy�����=@��áC��C�����y�g�}����*F�WO�9�@ݝg?GyF�?V��6�'��<1l��p%���-w�m¾L�`zJE籡P�s��-J�m��GO1���K��)�}��Ks�Ic!)!!���ϱ�2%B�).o���>#�.ss�������������A)M{>!��x���ŋ��#e9msm�^�|�q���rCܒ,D65o��U�/j��3K֪�����#����[�K��-}�ZRRҬcK5�\��H��/#�@�k���IlV�e�^��|�m�?����P1���:�lF���	�����f#�_�����!���",B<& X1K�v�q�:D%�H���_c���k���3<rD��;�~�'���Ғț�F16Ω߯�ۤ�ͻc�A�i����ۛ�n=�8ҊV/�CFj�ͭ?���쭼svvvsR�P�`��1	"|N�: ��e��F�ު�,�ݱ���,#cb���"�[��*���DWp�!�6��X��ᰠ�$����	JVWﾹ��O����ܫ�;7��[x'�����:�jg�h����t��{�lwsZbyM�>AUQ?�[P�X3L b��R,x-ūew�077����0��Ȅp*zJ�D�ƀ�>h��z����ק�I�	�n���!S�yb�R:���0h�k�������ODޓ�4��XrY6��\��CG�utn42t�1 �9tKQ'�$DR6�ě)'6�+a��P���|ۨ�!�>Sa�x����ˑ��Ղe�	ߜD����Ľ�l�%*�����7ʬ{�rss�̾\?��rz"<�_/��?���_�,A�����s~Ywm�H�=�@��>��+��4]��*///��#|��C�-��J<��L^b����1u���M�}v{{�	k#x�)@G�{����!�����C�U�w*�a�W"iUz�O��\�0�7m�n-ig���RLKK���3As�8���;"t��c������q�鵵�:5/�>���1۔F}���Q��\ ��J����7�� ��N��~P�%.���C\�H-���@	�a�5D�f咿��X��X�0q�ܼ<��s>�V������I����6�w��0 �oc�Q:���f;�)A�+�x����v�#9�Ҿ~�����XB��`Y굣
�J�P+��P5�i7;���H�a�P<��%�z�cbW��/iqf'^��=sGG��M��\�d�#Eb1Y㲶�n`"m!�O�7�2�L�	��m�T!��%Kb&br��H��7Q��@�yכֿ�s�����/�y����B�*�ڨ�=�=����'a��Uy�FD��!�]�����،-PV9�g�����?���׾����{�OKWg��ɨ��'��oeA��i��q�s\\\怄K��}�>}�O�u� �5��E�$b���ղv&��o� +�0̪%��#�T3/S ��K	]�o��־�k�Q1��?��tB�`���Y�V3�� ���u	��s����|�"vDR�A�.L�;S��e����%i��	��	��mmWD[����)�'��i86�X�L �T\\Ad���0o�ݛ��E�v�0�~�G�T�ײz�T��1խ��Y!�j��	�䛫 �*��M$N~�"9�:n�++
G�l�p�q�%���9��(� ���!��S�n��|r��[��%����I;{��k�kU���]U��7pܞLݚs�89��F��\�{�B�sbE&s��1��6�"彔��o|�C�6R<s���A�)��x�hkS�H���I)Zy�zp��/���(���o/�z�j!R˃ln�#�}i� pa��ip������,���5��4M�Xodm����Xc�������2��J:n����Oì	�$>���H�.�/��~f�<�h�	��yz��W���X�'�U;$�If�/7�$WԮ����D��^�X��35� (�g$�����~���s0������?-a0���Ce����IbCfN�Dą `����V��l�i2��(��P��7�ײ�d��^�Nb
B���o=����'�k-^�.�~� �1���(����/�|�Go?��4f�JJ��_ :��Bt��=Q��h
�.v5��x���i3c�D�gΨ���)]R!jᶪ��.^�����Z�O�Aī���!���#چ��|$vu��E�Jo���ƹ/k[x#���2�W�'�r���g��w&+��l�����7�+�x� j�f�v����F��`n A�r���q��>�5��Z�2it���75�bO��F�`e����m�o�p.H�-���;���it��ӳ苏8�K*��l���=+7'm^DR�<R�Q�r��L2���[�X�5�B��K�����{�T��B :"�2��+R�g�!q�7 �Ti�Y��K��X��o�g�~ϋg	�@f�w��`��/(k)��Ȃ�����-V�K�Ŝp;s���[^��1����?�^�t(�>W�Z�����]��v��,�Liy�'=�"�!��o��J�*��B���3��s�c��܍��*�YTBv-f�i�5��<���P�>����*oL�p���n�!D��>I�Q���u�򏣴n�4���6(u�� �]�����,~ʓ��� X��g=������@l͇݉ą��ݍTo
|Qo+n�+Ԙ��җH�:�}qO� ��� �&���!zΡ$��!�~U��!M�u��0>)�΍X��W	,u����������#oF�[�WR�9���!c
�mwH�B�!�}$}6�~T˕�1�����֊��ģ�4߫�������(ƙ���d3���Α �a_�r�T��_h�gl�d�ˋdY�/��9��,)�v�&k++㤓���i/hp:�W[�`�-c�=�}��l���W�:���]Re������U�)����H�ʁ�������E�� u.Нއ�j��g�{���d�o�4U�;0���M��8��o�~�$�	��"��f��D;&��l����V�ܠO�G:��Wl�|+�"�]湊����]�[��À��d�{}��������]��d�LQ�f)�	O��=V��%���@��C�	V���t)Y\Ta$�n(��D��Y5g�s�ٺ����W�)�xP��&�y���:kL^�ѩܩ�-}x�*��\�y	�5�m�.�O��5���# ����H�A�?�3�P���6�T��<��w�/�����"�0���{��&����M�Eڭ��3;T�auP�аKrl��s��*����5r���� ֭�8��n��`Y�(z���nmF�^ݮ�RNKN�Xs�T�I�C6�=�^ /��0¥7aH���[W��ia#巟א$�[��Ы�u��Jq4<W��+��%����b�z�!F����'��07'�,��+�M�m�|܅DD��&�
���-pk��e����6���l[[���\P@��n��٥B>��A�=?��[�����m�T1��9�yʬ�VϦ�͐��[��&>ֳ�b�GF��_�1[Ku�#�4<����^�s��6��f�?f��Lyrw;���@���X����߂����B������C���W�|�n�vqa	�:tmWV,R�����}1.~�X@�� \rܑU�pRH���}�#3>��.���H�����՚t��/$"f�@��vmMb������C����p���ĉqN������re��\���Jyx�}���+W#>C��N��]Ҏ�mQ�ø�pp�:��������gqL]z|<�R�ᥟK[�m�E�D�+�?����L���C{��?�|����&�Z��DKQ=�1
LY�Cm�xa���J�j��Y��]�O�n�Q�$�Rv����%y�����7���N}A09����k����e�(C��``ttt�~�=��u��7a�Hz#���|��īn�
wxe�Bc��V����%�J���Y�r�G���O��{CS��n?|~��xJD�7�H|����K,z�ﾮ���Y@c�s�]	��(J�����?E���/0�)�Gk������r����Jњ{���a�vRW�s��'�~{]�w8�X�-V�A +&���L���D^�����T%tk윲��u�Y|B|�:G��0h�l��Ǜ}��g�$?�sX���Y�w���٤�R���-�^;QhQ�I�X+]sH���;�%���w?b�]�ىq+�����ᝍ&���<:&&I�ﾾ�=C�������\�ܕ*V�8�����|���M!,%� ������`C�I�9��$Lq�	����ӵf��]������x��_Q�����^ �(��	��z�(tYO2�3Æ�>aA�����{��3U;���%�>�K|�>G����^s��} ̲t��6M�']�LI�w��E��n����m��ce1�Ye�̓��+���9�o�Ա�`u;��r�t��Kǐuj����9�K,��y0^p�IĢ�9�y���{y"�q'|���Z���y�=JѲK�>��٬��@|��=���
7=�\/0�N�PV�"��+�K� ��YA�?���buN��3xd(V��6<�[���;��?˲&���SS��VG=�=�1�1�@/�K��ic��揼Q�Q+0�] ��� p�m�-ƕ�Ǆ�U���|���7(��k�ŅzN���Sz�M�a%����2 N�[t�7�98�5�͏��6��w�#d��S�ĩ��:ӹ?�*V;ه�������&�D�|���U���%P���K���ާƻ3Юj�� O版O5���{�~X�x��2X�D#�2�~��	�vE����tq��T��={o���x0�ڠ�k�5�B?nHoo�5
A���� >ص��%���}x�'�(:e����ڡ�u�-�<:��.{���GmKq��q�)L���T��X��4#b���]�xX[I\�z�
7�k
��z��UF���.�)0�Ps���X� ���.����ڢR"�%���1b�p��<;7�뾅���9\h�kא�V�H���ӗ�ON��#+��s����x�l�AaZ"G�T�`�e�9a!�G��j��J�6�L(�8���/ *��9�yS���2���y�#�vvJ�
�kn�>S`Qn6��7�z�X�)�wq#l���铹T�?P��ag�.��"����襍/��<7���QB�sU�c<�l��	�����'��K��|��aW|ޢE��r�%ko�ç�6�v���b<r}~�`�3��ب1M�᷽)f����z�� 2o��H�b�i�#.@���
�K�~3tu?�5LA�H��Z��R}�&b���$�x�_��ym����C,��GQ��ߦ��
:�Sݸ�J}�������l�=6���0)������I']s�W*��#g�pffwP }��͖M	�w-Y�gm�(�y��E%����aҪ]��,��P�܎y�p�m�����nT��ܚ�|/�)jI� 쎍�'{v������Åg=�x&֬>�g�W�*�L���>k*��6�:�v�O�FR�t3Ͻ�P.U|vb�����*4�l_*�lY�͋��2�i�+&\�ܵ����C����.lL�[7��5�F�dBd��mc�����}������}Z���t$���6�|E�����F$��ːQ���nF8z
X��M� �u���t�텭�����?��cr��� �wA	�S��Sl�.*.�Us5����uB�1�0<-������х@��,PA�0c	�y��X��e
�o]���q�Rˑ�_��o7�t��ɝXL7�ԋ�c~C���U����7S�/�y���G�zC2}Ė����1��F����rY��*4Vx����f�W���ɻ;���0�>CW���p;��q"�鱏�> �p�?|i���K���7�]sz�'\3�;
y_X[Y�鰿6�)ْ�����@������0V��"Pq�Iq�9�SY,��a�c��y�n���%~{�*�6%����Ju�1d��D���Q��B�\Zc	v���7Su ��J�&��b�������Ү1r��t�Bi���yMb���n�e�@�Q�	�}N��u�Pq�`Zi�v�.�����<����3K4����P'S�Y���s
�h�cA~L�]�|0���Hv�:y#��ȋ�까J�Vt�X��	zy=�Ų���=?��rǵm&�o��-��g���a��~3��� �q_u"6�}M����"ĺ�ǡ�|�1�T)����sA�DV��(�,Xʒ� 3o1�v��u��̾�o���.	3�ih�_b�X �}'�>C����8d4�9�Яzn�0/���A��'�����H�Gi{3�V�����8n�0�kY$?4b����
�n��0#�J_���h���O���Z�\ �r��i��<�Q/��[��&��-���}��
�J*�1m�E2@���/>��A-ၝ�Z���|�����i_�o��Xd��f9�]����d/��%�s���Cq%�7��R^����U<�ؙ�4R3cP���)%��}���I�!z����q{��~�뗩�⢈���\[	�~���C����@�x`�aZ���.�l-4��q���J�B���ujӘX�˦�8���(y����n��j�Κ�ʷ�<0&k5��%�yQ0�0<��B�)����������^�E�`��<�0�+�3�i���!;F&���
JQqI���7X�@������]"WS��R��O?V]�b�g h�������/�w~�.R�w/�P#�l)��>�{��َ�U�Q���l�PMd/gv��7rlؗ.����<<i��Ծ����+9��l�]�L ���>�S�g��T��/�ow� �� xoz��}��75�rq靤����J��ʀ��w>u֘���v�t3�V�`v�KSR��!�Xシ�n�*X���I����g�g	�5 �� xc�ɚ�嬥��x�*��s��V���	�����f�3�l��ᚁ �F�y)���h���n�����B~{��Sm��jť���\ e���"�v����Y���mAp�t	��;o~���W_�����׺��#&+Lm ~�6=�'6�����,_��ƯRe�;@�ʆ �v�? w�)p�ջ~�Q�M���t���<�(����)]���~�=��\v�u�9�cS�nD`M�QI��1dn�������b�`8�K�z;s��T�qR<,����u���*���XAL���{<!�;9�%�x�L������*�?�¡op��Ө�~���J]�e|�e|m���b\�$c�3�;���'����`LdE�kY�K�e����̂�O�˹��y��d����O�!e�HaH�9�	�A��~n-T6%ںhR�B|�Ǘ7��U�8�FmX�;6~���8�3���i�ha��(]`�/_�}�K�`�=�J�@ǔ�촾�6[z)�}²�~�aG�@��j�DT#��1~y��r�W3�ꏰ����R5㝗C���Z7�8&+��0�� �MF��8U8���c�F��'�Y��W�=\SK��{.n�Rfu��%Y5Me�s
#!A��!�6 ��qh+���V�gG��}������ޖ�RTS�ڏ�J	�ʋ�\�EC��y��R/���q�-U2.��LRn�&&Se�b�E��7D��-տ���X�І`%�{k?�{��O4<��Z�4���>�vC45�>ʱ��%o������ݻ'����M%#��.+n�n�E��;��w_�rB�/����7)����~n�B�ou4pF�{�t\9���.����]f+�h�����RZ�5/Vӆ�m�OW8��M�nf<��k]_̋i��4j�]�\��U����/ar[�OB��訂���뀭P���]D�m��H�^�����>5�:*�[v*�%��p���,��GyJf�iiz�:,:ʾD�"wk�|"�:���p��8��E#q�-V�q���D�&�fy��f�g�i�$)a�z�m�B��`�O�mˌ�x���e��m�J�@��t�/=�-�s�U]�:yi9~H���đF}���ub��o�LԞ��v�٘�
JO��Y�|�	�)��p�=ט�Ղu�q���+��{X�F�Q��i���� *�v�[��\�ck�J�l
:�w}��s��y+YNM/���ќ_[�mJ�2ժ�Q��ɾO^᱉�%�>R)��*�=ʫ�x��n���V��
��0�sw�7mx  -2([�N���SpqqiN��Ϫ�!�ok�.E�����y����0��eS�ϱŨ��p�:�4���7b6��(�?Y;����[zq�L.��5B|h)c�=Wgёˊ��ɆX�n+SUFaa�r�{(tI�r�0�3��ӞW�lD��q��D#V[���sX]�=+Uґ�Tu���?�uȲ�:+̈́�\ʻ���f�>�T��{��t�,�.B�J���iS��;����e�$�) H� �z�HME�
Y�.�C(m믏��=��>�_�.�
Z��>笞�!��*��ZO�pr�+Lē� q��	�FN���|\���nT�x��Sݱ"��lJ)���(�()5��+��q�hM:�r2���^G��D.�@��ʕ+����K�;_8:�R\�^){[9��/�0��y�e�:a�挧�������6��c�Șr,s,�� �ty{�\t��Da�����V	X�~R�	��C�������ue���`!!a���M.�GV����/T5E֨�t4� br%��R����,�໊R�wnp���(p�>s�Pk�$]��>=�o������*�<�0���6R��a,O�+�YU��:2S(�Yo����Ou���j���٩�*瀞ZXȫ[dڐ�K"�d�Ф���q��G�H8tG:�
�T����\|A5�BMDr�꽬���������\\���QQI���C�ȩ�=2)LRh87C9Ξ�=p��f�^��$��}Z: ^���>��F?}t���������ze�D�+�x�:��������ӧk3n��Q�~5Ō�BBB-o)��W�[i�B�����2��O]��`��T�$*iVDS���e��wsu;SQQaҐ�w��J�, :��Q8�[}����Y���?������B��]s2[3A��V�4�I�{���i<�S\�Rw�@��S��Mz�����ީ�l�8s�n���RN�.�b����̖�ȹ����}�S�}a�nCm?z3�'�b��C����!3>�K�������������nnnT44�YK@����(<���vh}8PB�SNIF�=v��(�;U-��)t%7��|�>�����T���&����q'����q_��mz�}����&�4�o��e�.ZƗv'��S��YRM��5?��C~ւ��=��P�q��-��8�%9
�#�a�����	^��Y(��8�����
ϥ8�Ja׺�t�� �!�Ps�?����'�-�#:Ԟ
�[ƷZ&�6�vW������ե{�h6LW�UI٬ekhL���9���"��mu2%99���)�.�(��q�'����� ��s���jj�j8��{=D��gHد$Q)j �v�����G�Frjj|e*nЪ�Ewv�UzB��0^����?0��C�@�^W��qwp�H(�49�`�����A�ޘf�\�H��b�֜�̱�F�z��H7+ΩꖆgK�y�Q���W;C�UL���c��"��ȉE	L��U
pf��4� ������sV(���N�揑���ǚ�r�M�#�G��YRԏ��|�W��%o߷9J̗��"���Lֶ�m�ST#���x�;�4�
����� �r�MʱݩѸ�g�SeT?���/$�wЯ���ِ0�[M�f+�*+4�DB/��C���z��ꠣ�a����d�����l/��W5�E�}wz��d�~��AJO��ً?��W��$���h�\Rf�Ђ/�m�|�k��s�E5�я���5���!K��-B���l�
��񧅖.ԧ�>,�k�Ύp�ė|��������3�I�Ӑ����|\�/Xic8�����'_������T�Ӓ[�E(m�X� �Ӽ$�(4��QͲ�����Ix��S�(�M\~����k�K�,���\���ݗ)$6�� �
�p|H)q����n��c�b�|��&;��ܻa�K��_y�/̩P�?M�ĸ��5p{��k�,�A/1*>����|��It���vh�M�_��S�{�2}�	s��'nN��95����Œ��c�|Ww>rQ��S���{y2�=��b&��W����_��r�<���8�NF>���b�>�յ�=Z�:o]�B�[�A�4J��L���՝�Czzt�D&���$R-U������������2'�~��Y�-;>W��M�������Z�O帩��+�#�Cj�y�q%�!���>��3��s��+A�=�9���\��K�@���8"��՝ e�΃��=V�up����ѳ�r񜨙㩆����ґ���V��Q~o�P����fle��4���	=}jX�*#Ø#�XRÏ�,���lFMXnou�,�Ki���[L��p��=l��j����ל�$j=P9^�R��覽13f555�+�ڛ�)���::nvW".����()u� ���
�ni���	�Ô�?>���t��]W-֐O�ޙ�p���s��e���%�F�<u-V��;�
R1�'�q�ᆯύ�ZL�t�a%�lg�h
��i�.�h��Q��џ�П(z��������%�1o���@�r���z�H?�]cz�m��GF=���$�Y���_L����XE&�#Vr��~G�ܹ�ǒ��U&�a_��[|!C˛"#O�����c�7�4 ?d렗g��QMGm
�E��#�t��7�^��V0�0���7��;avB��$(8h>�v�e�����Gx2�i>��ƞ�ta�'O�:)f��o�;��������~B`M����x���͕r&Z\�2�*_��ڌ�I��œ��9�a,��;�9��87�82�ѠW���*lҐa�+��zЛҾ��XU^L�?���Ak��n����\cv�&���zn^�li)u�r9��h�l���|nYaPZZ��<̈́����AM���#���a_=v|�+�(��k��Ž�Gx	��S��>��b�8�6��e !�D��� ����rμ|yW�.<]s����F�q��N
Vf�f�hֵ	�qVJfN<x��ėT���L^֕��Y��&��s�h��*�r{�-�殟��]7{q��1��i��XJ3�+�`�;�8w�2�|��ի�U[I_�S�tP=Ar��AK��K5���3�6�k�V/U����d凵EH�#�qϗ��ئD�X��v�A�8|���oܖ��gs��3$��ݱ�"���`�$!�{q�`������ͤeL1������y8>��"QF窝��$.A�o!�� +�:��nx�{+N˱
 &��81��O#3G_D��%��o���ߵC���$�@�ab.)�C�fc�����G�],j�Y�tw�B�����
]6��օON�[GAW�u��
8m_�ui�ŉ@�Z�����MǠ���a��|�	��_!vfSg�V�:w5̱ndLs��>��a�tyb9Y��%�%��o>���
nte��l��\,^��ؖ�豮�lPGṣ��ݠ3z�;o��|G���C�Z���y�X����<u�nX2ܝ('Yf��L��Կ���g�s%�s#����h�6F�i���E�{�Ɯ���� -o�!�v24��Q�;X*&��n�Ǽ��G��Of�I@��@1������9�M&���j$��ǻګ֌�'��Q������k�� ����TX�8,\��S(�,�Cա����o�Y�N��]�_���vUm�r�7*�_a��d,T^�G�gM U@Hsmkn���=�C�X*��AG�����"�h���сe�N��B�����Ɇ�?iCV(k����|�I�� ��X�Y����d��)�����mi��+Eӽ�=�� �=ڮ�F�����h�}6@c��r�AS)t��z#���h0�ݡN��|6�syȣ2x��gd�0LTr�)5��������K�	H�mg�J���s�,�p��Fc
�Wɲm�Ɵ)��om�"zCY��!�֋�;.;�a�.cR�X%t���e�]]�}�m��ZV�q��W|;5����9���1����J���x�;x���೙Tڟ�ԕ�Z��dG�0j��"x��A�=G4�.x�G]�Zżc��T`ӆ3ޒm|�������ug>\[mҭ�s5V���j���ԡݒ5��҈���9矷i��s�S�K� �0�NL�7f��В��B��]Ug��)6��gg���LpM=CJ��hT~�#�VG�m��X�S�!�H���
jˋ"�{�5VhM�8�l��w���j�������|��R������o���~z���[쮍s��`�C���%��Bf��P?�y���W`�5�;����c[�lf� 0b��p���Qfc�/)$�ä���B�$���fi��uS��gu��X�7׾�ϑ�x��z��E�}�����Դ�;V������C����u�"C�V*E���.ƞ4L�|�Á�[^�5#�S�m�=���l1�CɖL�.TRW~�^]R7�_��pr�g9�_.��M�K��H�>���N��R.<����hC,�c�G�4�AN� �mpii&q�'�܏%�j�	b�TTx�[M�MoDa5�f}�W*���IP����l����q��<��e���d��$�=yo�%��<D�'PX�d��&̋$���`�J��ﶔ�6���߉g3>�v�P����٨n���;��NVF"Q���ƏCʇ"����'h�藺+K!֪��s����	�{��]шJ����#7DL���ǃ��s
3&���%�|8U�<��r��Y��ܑ8��}�u0&��N��ܽ�I5{�)��[����y�4S6��[5IL��u�:h�N�.yg��NÍ��_4� t)����d��N���z�vq�d�����r<Nj��D0�h<�ӹx��Z�mF�D>�!���ق���0�6D����{���?rhFW�����4̣�e�'Gl��`��czoj�u��J���C�5ߵ�?�Ŝ��>N*�����Hy5�u�N�*u�jn���]y�ēD �����������i�)��T�[�%�� )*�g�轓SR��"i�>�4�Ј��[]�Qҵv����æ`"���B�2Yl���J��9b��%w�E��S�tJ�����=��6@Q]]}2�	��&���yA?0��3 1킌}˺�2U�X����sA%�t��)wy�֣@G�J�ab���/皨2,��u�L]62��.�M��k��{�Ez>�#��5Ţ6,��sL�cR�WQ3�]@�a)��[)L��*�z�z?zn�7�e�8)Êsk��S\l�!��f�m ��m
����Ņ�������(T��ɗ��78<��ì8��
��Au�q�8��tM�ϖ���|�Թ�>q����x���?��4�mZ���K̨�۴rz�������&��Y��O�D��4�<�'�8�Mf<H�҂�dvVt���w�pQ_���j�-h�[��s��f���]x����N+���rE������*�rc����t@ca���SLB�{B�zt��̡��ޤ	j�.\>7�,<����;��k眗 ��k��m?ǎ���&�b|p��';���՝E��Bn��*�%rZ�Z�Ň�ǐ�1����60����~m���5qZ�w��=J�x����ّ.]$�/Ƃpv��vϟ*ph|h�ܧ,�o�K��A�I��"E?� �v,�G��8��#>EDP���b���ʋp�D��9V�7<k��	SU�>4��dLAEb�Y���Q�`�����OBr GI��|)�[���Eu��R�<���f���#����ѵ�(�i�b���9�K
��sٱ3���f�۞�����lw�yl�֔xϯIVV�F����o�B�;��:ӑ�싫\C������j�Ƥ���椱��\���!໔�	*����rd��{ţ���e�'MV�v��E�s�z�� ��6)�๬�kI���PY���̜e����[#Q�^r��'�m�:�Mf%�1��G�E�� Z���;F�̂�S"ѽw˚���5����}�Bܸq�sG�
S1�m�����Eノ���@����$� C�-����$�sxX� +�}:��u�2���W>�9j�����t�u�U�օ�%y`���������5*�g�Z~`��������� �^갏W������3e��9`5�I2T, �Yv쾚 `�0��BC�����IQbb��0����h�-��|�o��Md�[6�Z��N�RXҪ>�[��D{cZM���������+���ÚC�l@J1���"Lp~<�n���%j_�e�z��쟎=(�dyl���ȼCR��� ���)�K�Q6�����>�$�{�����Ǆ^u�Z�e?��� �n_kى2	΋g9+�Db�˿�~���_��q��'���fk�>&$�O����y�s��p��6�ym_�����gvR�-���q���q��Ecm��8���Y�H�C"�a
�r)��M�X�n�'�Sn}�U�FN��+�ܛ��~���l��EX1�F��k`�i����3
O~��o=��q��	��I+�KI>v�4V���L��BK���=�[�wcE���*O�����T����bF�L�A"�dgHlI�
�h��0U\�j	�:�:�[�ob���G���S[ ��k��8�>���T����`A��=�%���_#��y"��{�ԧ�����D0߯�>ԣf;o��
y�xs�,].]�J�O�m��|R)�kl!��� ��<����3^\\��h_�Wl����]"��+��@������lоC�I_��ru��j���	�|7��`�ӛ���-V3+KRSouvu��T�4(����b�X#�r�j0�h������]]0M󷐗�F���wd(������yX�҇�D7�Lm%Àژ�D���G&| ��R��Ϋ����xx��L"�S$��0���B,�R >�z~e6m,���ur~N]�]�m����*�صԓ`_����12::+)!?a�ʁ*���AC���;}���W�[��wԆ��Wu�����U��p�xǲJB�{�[��^�~��A3?���ԋQcF�F:Uo�j����3Q3���#�h���FW0f�RU��I}�A��^i!�
-���[SHm^l���J�TW[caDn��}��8��1	4fR�yQ��1-o���*R���Y �wh�k7s�D�r6tT�O�o;S��ѹ�b�D��,wh#�m4�u�m��N<|�>�I7�O�ȡ���z/���1M��\6���s^i�ăI%!��37n��I�%v���f�4Ynk+���i��h�D��V�so�g��4+r^jI�F�DSG<��۞���?.غ���M��o�}O��k���VU�1z9��یwn`_��]W��D�ɑ-ؠQ�Dwй����F���@@��.#-�N#.��dv�А_e�	!X��Yt!ܙ���^��4!��~��#k�~T��]/@^��y� �g��Ւjr~��,����N2��n�jɾ��焚��X$�)�`n_U�x��釟cW���˽��j4:7w�ٟ�a9�%�P2B=;Ce!y�9o�>;ʿ�H�����ܑMQx�F�v
)i�u?�?f�^�_�4���e�5<�m>�a�ZHd�0�E�U,
�ؤ�-���Դ�݃Cc�5��Di�j  �j+u�J˯�ҩ�o(�G�;��U���FU(w����sa�_P��_&��sI��څ��F-�� �B�=�S�Hj���<�￹*��u�������?{�w�ֿmT���_��j�[1���<�)0�F��A����+�T������i��I�vz�g
T�3����>@�b�r5'���j��i���5E���#P����R�s����������Y�T��C!)�풇��?��gXS��7|EF, Hǂ H��q�&]����;fQ�
ҫ"M��NP��{'	���Cy�v��?Ɠ���������]�����MQ�s��Y�a��@�L�䨿��������!�n�
��E��T����� �PK�t���'p�ۅ�c��t�~ <�i����`�qd��(V��G�X��q�t���Z>�xp3M"����U	��)c�0m��qm��wWS���ܩ�N-Yoj�j���������g��?x��	���tU��چ�}����T�?4�O�W�Xw1F]��IY2L�W%_����q�7 �ם7 �8�A[�	à��s&[����6��U�>&�(����Hp��d��L�fW��e�co�n��h[k$6�~-���H)$���]S�/�����ӝq^ɑn*蛁2X|�`�d�{t��f���?�י��Vw]z8ts�i�/��7������̼����������U�?�赊%kfJ^__7��0���;)�y�Q����sf0�:a�{�]�?ə�[d͝�S2�]�݊L�9��]��˧!H��Cߠ��o�N��pY����Y~��y1#Z::�{p�?��=%M�:ːW~�*����/6�����W��@��d�����bR?�]�-�:==-���)����Z|�f?�d
v撂�=�Acw��T��q�'?}���<�@7�}�����URN��6��n$��8c��E����+��=�˹;F�a�1ێ`�^.�g��ny�:��	� y(��W��Q������ZXX���g�#��������X������WN��o���q�L<xy�C�"׵�w����P�+wZ������?���Z<����z��*ɝ�{ֱfKW[[�/�s���y�qOK#�/O6��v��e��Aq�Ax�rg��ZQ��D��bֆ�5���[�Þ�|=װ�Y�6��ɟ��_Ϭ������bv~hC=B�����g���gn+#�a�y���	9�
.�m%댻�"%�Q5^[��4ڣ�v?n�;�e:�|�>�W�,h?LW�}M���������(��r���ݻwѣ�T>აQ���5��lK��n�ܝ^ `kr���un爣�7B�������E��5ɫ�3�彛���#�T\��"�N��^��{Ù��D"U/��!��������j��LK$��'߮b�|��U8�q��6�̦��-7�L��\\\���+�em���l�z}C8�Ib��/ ����+B�����36��+s0��/�fh֌�i��+��s�8���<1��ϼ����[�g��7M�-�9�ܲ�7g�Hʨ�q7��P󱴴��v��H�R\�;[�"���L��n�1�h�6��FPc%���y�S#��\�[Ȫ�{+E��~C6�׊^�T����vÔ���cBJ4��bU���&��]a(������憂��~��%�WK�O��}��>�'�KB�<�Q5�Gx����X�O��nmp���G���D������#�C�KߴE�e1v�5��p�:���+���	���l;��Բm��ܘ+fE}<�joƻ�~�޸ULn�?�J!�7����׋Q���ޗ��᠓ɩm$��0���I�wU6�Hn��@o��t��АT
6���q�u$~���ѐ�ɞ�"}Xm�����\p�z�M؄��b��{b��pU�?��#ˉNL&�i�zs�O��J/��ܖ`�ِ�O�'��ΠZ��*]9�/2,�5�T��Ν;��}.p;�|Qxe)ǫ�	RSH�L􍫂gN�`力.�"yk�f��.����wM3��A�UDb{��t�d)�Y��7n���#T�(��N/���W�F�&�ô��jA��EF�����wWF�/�y�D�'�}}��r����O�ݻ>�q�])�����O/�c&��o߾��O;OJ� �{^�0�gj���<�HO�d�)A�ӫNw�9O� ���P����#�G�X�g9���uڸ���Aq�A�m[��_(]�ٕ%z�ș�bVF�Lʀ��MvD����J��B���%�p��1c{_is[��-7S�02˦�PA��Y�4
}H��㦡��`n�RR-ߪ�~טQ�Xyzu���S�p ��S������M4�s���	s��ѹҠ�_i���)
�0L��J�W��qmv�r��\Cz���\�˝e5�p?��T��e�ꍜ�LS=\��sI`@�6�}/4}���v�^}6
��CbY444�����BBoT��P���U��H䶰R#�	P�R��|�/ݵG�/�����V����H#�.��'Mw��-��pP���6w�}�ٶ؟]&��Z&��g�pJvw�m��-U����iҶ_	�P��j$��iMo�o���ʖ�Ni{�Q44�*��l�j?:��;�>Qc����:Cds�^��<jl��,�ZTa|�t�$���L2@QmLE�vԿ;��*�3��_\�/c	<Yy�+�}�+����C~���D�T�'N���,���bvC/��R��Fk�Y�x�^�측�Fw��b�F�K-3V���z��3`+DП�=�Q��&/��U�Mxy<Kd�q�jz�I�p��0=D�SRY?�K|o|d���?��j�J���N���b���I�п��9�F�̟8��1�����0����eb�b��d�Hg�,����� ��K?`�������`�6�� S1�'���/��x�����@���Y���㴢o�Ѣ1�V		�Q�"�h���~����z�q	g��%�&�҉}˰����$���+Rׄu<MD��!�6X���BUIA�������?�I4CڥW-�����_l�J��xO��e�ʪ��_ۍcMO�ŕ���L�#'��\Ԫ�>R^݉v�l�0~&�|Ʊ%9�ַ�Z'cj���u���n��4+���J8[i��?y��ɤ���N��n��l�c�娅;qF�{[Щ4BT����|d�S�Ў��$����l�G�ͯ��X�&2��d�R�=xY��s�	��n����%O��Hc�䇛�g*���B�Շ^ ��5ه6���N7��W}1&�N�G�tT�D�������E��_:{�C:]�ZY%V��[7G��!W��~��H���+��s��<�,�����H[A�jG���]�����y6�+=��_����Ք���^�0�5<)bSW��Uv���rcF��%�+Ȳ�����r�={�������-�9��O��E�'u���,��a�:O��b�K����%f$B
jd
�N.?�������_��ˏ��S�*B�v]�3ڳ�����k�G/%����'XX:�V�Ϗ�Z�\T[�wh��^�87c��(�3�&��+Zg\�Z�J�X�A-��@l�-m�	ſ:�߅�5��5֨�3��+
��4.�&j?�{���v:�;�0��_��J�o��*��e�Л��i�:�Ä�%���oU���y�Uصsk4��|���V00��P��*T+q)�2��n�y��D40V���ڽ
�=��*c* ���ߕ�1�eA���Z�d!M5U��r"�P&H��YE������B�{��rJ�u�����p]/�o�o��5���Vc0���5��V��HTM�k�EQ'�'��F)�gO͇�9f���],:��\������Ogъ���'Rv{���\fa[�+�����eȢSȄ�O����Xn�r�4:���%B���T�1��t��B���A7W����Ӌ����cj��C^_f���*��p����1%�@E��Ԧ-Æ���~)h���o?x���\��~��^+ n!���[ث��iUN�FI�m��M�
F�u�u�*����Һ^����#���ݥ�ZQ��=�N�f��?s���x����������>��vP�F�n����vkD��5�ӅЭ
�x��;Օ�7c���S�J���/uʠ�N̔`�*+_�(w'�4�|J��US���V&[)�Â�T��)IF����H��w�a�M�9n�t�DC�I<w&m,�eׁF�� ���	�2A��.��.]��n�j�9��
����ͩW2$��x�����؛�.�gq��o���$��V��Q
${;g*�q�3��$Y�6G���b[V��!��ԃ�� 't�7�wa�[�̶��-U{�ZV��w����l|�%�g_	re 0M�q��bW@�y�19T�P ��q��%/riL�Nڊо9�qg���[M�]�3���"	��W�c�m4[v;�@PK��-F>Pz3j�4� 1�����"Y"�t @�� mTG�7H� ��s3eisI�}zQ���^�
ڐӳ��a�3�qa�b��V�����75_�m֟�ON�/��n�u��^��V�h�R�v�&���$��tf������R�X�	M�00�?!͹'����!��#>����p�>��p+�LO�ן�ɮ"�,^9���k�ra���3����ֵ�nkC^���3ˬ��)� *~�i�
IݮN�p���¤�I>��(���B�j��,�E�M4X5P���Kش�E���ӷ�:�;�8U�)��)mw��s��_}��:�n5K�A�{��,�$��z�A�?�6uƐ��hY:B*�;�_�O�n�m�� ���Y���WՀ^���;�U�.��Q�o�L-8\	KHtʸ��t���d�B¯s ��̪��	��Ze tƩ�$���Z c��yHRdɐ���/cǊ����+Ɂj����.�G�}	�����}��ص	Ξ3�ޟ8�ݦNVV�d�B��̊�K��笗m<� vNi$CJ�ތ`�"��A�L�z�n�L6���_��-��yb�b[��@R!�D!�������N�iI�qY�o^�]MM�&��1B�ܕ	S����K��`�D@Q.��I�"�9n�5��VJn/�Jb+$L^�n=GO�(���eT�s���S��or;������jv�z?	�?e����� B>�艍�MXƠU�G�k\�ՊV��Bڮ�b�P`i��SK�y��v����~�;��Ʋ����~�\�m]�97#`��c�%��}�u��	u�F����f�[wZ/��W#9�W����xz���r�S.r&	rrrBje#@+N�Y��%�?� ����K���0L~z�V�!'�T�"��toXR�8/�9��Oa����H'S��_V;@6��T۬�V�Q7���t�"�:fp.u���._茇o�Ɣ�����n�,	�B�#��E�U׃�
߸�l�񽒜��3﹯��
���.q6���KW|u4~�_Q�?$����]`����:�Pς��;����a��B|�X��,��O��s"ތ���?%In洇?����OpE^v���1�+n��	1G��l^�6@����g�υ���et�Cvr�*bТ�S�j,�!�s�j&kޑ���3�k ��L��ZU����H�u�.5�I�1�P� ��e��h�������ϡ-T<��7���s.X����~,�Dw�d)�|���6}�כ�$���uk��Ҟ���X�ʲ�$h�Hx	�҉ JC�ъjjnʜ�IXt�Ĉz��a ���>3���{=[���)�h�Zۃ��I���
���
�ޫ���s+�nA����J�lja�r1^{��o�˗`[�q��E=�1k�{F�ZHO���Q��s���Ak��U���sM��{j &��,��ĭ��(a]� གྷ�Z���}��OY����S�8NԬ�����R��T/����k�
T�ɒ�W�j+|��k�v������W[�z��z|Ǟ�R���;�ށG���Sf�' 	���ِ�ʇ��<&$wXD�d�v�*�z��id�R;�����y���-�G]�Ɏ��t%[��&���6�K s��j�v�է�GgńQvU3��3��e/M��/D��yFw����۔�c�M�n3�Vg�٣��S�2����'��Z�/0��.�IO��р�$;�_[������հ��]����F*6=�&��E;rU-1�F�[�W�A[��j�~ޠw-4�q�� �gWW��N�aT���Ql�6L����H^Y���ȹ�V��`�S������W�(���yR)XVdX�R���}3/�G�((Ft�s�;�ա��{�e�E&-T�Ɯΰ�zf3��U���;������U�5���?,����܍-�v��G���y�|�q���w�4=�"��
; ] ��d��ОS<;��wWG����K�Ә-?�����e��D�#O�f�3��CT���@�$LvW���:d�N&���������>c�>~A��74�'�`�N���{��|)�9D��gn�D�v�I����a����HX���5���h�DT�F��A*���p���� �8�8��_����P5(����U���K��G��o��[�>x��8J���flc�/�2�Jne�8�r�^�5e��*_��Du�g'�s��ŏ"[���\o/w?S�T �-~XQ@B�������!au`�ps*�Q�D����X�,���8�w�g_"�3I,��>&��4҈;�C��1_���*�B�ؘ2;���)-��=�HD@�6G���cB|��.=��?��B�8����>h�b�
�|�3�>���7fcjm�z�/4���㗤s+�ݲ���dBm���s�=;~��W埠�y����m͖T�<L�_N��7+��vЎ|�:���]+�E/t,k�a����>"w��|jL��I,�r k�?��$�0n���-"��`��4Qz�w"W��\zs�&��c�KHH�&]�&Y�/���HZ�	:w�Ŕx�V̇x8c�1�zN[����#F+��zE�5<�o� �i�m���m^?u&��8a�%��FQ-�)����NrC �M�B����Zu枥�v��_�!�P�(�a�7k�7nf����d����^)	���
3��*�W�Q����a����
"�q$A�.��~�WU��td�z�'�l� �y�U|�a�>�����Mp媧�C]�Vb\)��Υ�����P��`t8׋��=a��8���F�x1�������o�LZd'�é#i���қTYۛoľ���%yԉjI�Z(�����`M)oV0[e j�o�Gjq��<L~�/TC�N ��Ԗ0�ݴH��r�7�l�D}e�k�1l��K� %���!f6N���k~�i��9�����ˀ��� ��I:F�
�6�ƺ�9�lX���P����~3��YE�3m�]A�^���`Vv��W+z����'�������ͭ����N��v���}W��>�O����G.�P�ao�p�{_��^o��@���D{Ƥ�ki�Qe���惪6�]$���ЏU'ǭ�)Ab�:�Z�����|�zt�����S�����2�uCVd��<5>�SjF���^�K�����D.�Mi"�&rB��4PuN��K��W�q�` ���H񒻐��X�?x���-Z��Xc^M�u�@j�A�W;CCe�2��g�7H�9���gW�_P�B����]�44��'o��~V��8���9�e����}�0�B�㠗�+|כ�13Gj�Y�$W�}�p���Д�Y{����^�
�j	���v�eBg�_����Y$}3�ؿ�઼]Z���C�S�#��n��͆�s���a��l�Ķ����� 7�.θ�j�%�"@njP�	fr�ns:"�%zC�s�����jIZ����^�֘����'��m�z���S��2�q��%���2���F��'gZ��S��A嘏�wc� ��v#>����A�.̖�S�Qn�t�Q#��<�����t:�N�VhV
��mX���j=˫b�a�}����p�M��|�L9���s����%kf�F�{�*�����V6�t��1;���p�H��X|C����l��I�%���u�r����:��Sh�|�Jn_���{�}��eB7fL`"$bGZLj,�J���yrw�o��e�W�K,��r�~ۮ�0{��g������VMdd�Űz}��f�
%f#�y���ȅ�LճIǎ/z>��Cc[}b����)�U8�����6���F@S�[.\�OƂ��&����Gb5tM��v�ʲb��۬���Z�i�)e���ug�ACBx�	P�?���OMu|V[p��;ɨ��դ{)�&�1�6N`c0�Nj[��[���5�>��]�X�X��l�Ns�+����;�����U�I�*�O�����;"��;�AyѮ��7��V���b�G�A�� �F]\���}��J�s��`}��H?&���2Ȏ.��]�t�َluEd� ��k�t#5#�g%�� �����:�:1��
0E~t͝�N�L���`è8!�j�� �2�"�v��O�Mp>�vI���`���)��#����5��00�kw�{ht$�?�\��Z?O<�9����c�=��Z��9ʑ�홴�m�%�j1l����L�15�´(�[�CwK/���J��Y�UKZ����F���;�2�L;�֋n� ުA��I�3�Iw�������tu�e]��B�w�g�
9�:�H��lѼ��U��ɧ���ϩ��y��럪?��OZ�{�R\�Oq�t�꽠��n&}}6@�e��Nj(��v��B>��LRK� K�[��5�_�^��.�I�E��#j$���W���l����O��)���WɆ�l��
S�����>��_�{+#X�X`��p��,�u�u��)ޕ-�؉���Jg���o���r^�k��e�ο�Vyby�]�j� kQ6�}�[��9���d����ԊcĆ]��}w^1?{7�}����,c6��`'�P�Q4#أVu26vl S�-*$^�S��'`���c�m燧��y��Ђ����������G,���=Y8V��?Փ��/1ozQ��l�5�G�^L��&~-ɤ��#>��V���n$}Ό��=�৿�T.�g6 �c`)��b�(qxXg�1+E�K��6�E0pTB�W.Y���7A3�{�L��aa�
��9躵0�S>i8�M";V�#�t��CK�շ=��f�ӟuP�S�r�=����7A�������s�fP�)�<��M�x��7@�ط��eF�s�g��@	L;�4�Za�N4\�<F�(�+���W&�voMd0��hX�H�F�lٖ?h$Ȉ��j_��#�������L���Ͼ��ghⷁA�O�,�)p��e�lv��e�M�IT������Q�8I��6niG�h���j�`E�ט��B�B�� �?�3e��{�k�����ì����|��F{�I��a�`_q���U_�;��Џ���������K�xg�^��! V�U²�T�F��*�"WY۹6��#)��32�l���=-#���no��j���W�g8X}L�h�n.�؟�!p������Y>��W?;ҞX����W��r]�~�K-��'������U� ݀�����c��*�Q���������DMy͸J8���2�\�,���=��ZS�� �?����B0'�5����r�+�X�Yd1�ܼ�w�V�[�j��=Y.m	ׅj���C�@u4�wbL�%��OL%�NA�UJ+���� Rz�1yx�������/f�2��,{?��lw�\b2qt�K{Aa�u}�c)$��U��P�iI4�6F9�������H���sKz�ʶ&��5�TB�VR>rdG	���f��w��SVy�-�U/��\}��_��Zl7V(�P�i_�0��J�����k^#{�S��e�@�yGۿ���L�-�̄ĶT���a�HP�ip����hZ�EO��	"N�S��ٞ���Rwr��g���ʹ�͚���%�5V,i�ԙw^�2/p:��/;paǻ�Q�������m���ۅ��+ hp]��,��ov�� h���or��(�0��ON���}��^�3A#�w�}�ޏ���u �|S�d���%��=���R��(���|�V��y�qN�,����ν�Zz4<�ϣ���r��b�����Ƭ��{V�� @<R�	ҫC�F����Z?�7�0O�״d�^?���Vc?fE
�"W9�X�奕=P����C[6j�I�*�$o��}F ���=(�Xۿ�a2�^+U�^s+�7P��S��w�;����W�0L��V��Bu�x�|�b���c2�\&�^�w���}^�,u/4��3�;K~��M=�$̱���U>pS�+v{6XAl�4�� ������0���:nM�@�X�5Z���ȹ��=O���n��[\ZB��5���3�ɺ�W����7�n8�BQ���AGbd�������SC4�9�3~��[N�tX]]��e��H�� �&�YY����$8=�fZ��_6��l�Ĝ��C����;-n7�yJ�N���sy��p�\8�N���G�G���Q�2��]�Iu>���}�١X�p��c�ܠ�����L��R����R�7�߼%���M���'�C_��9��'f���XL�~#Ʃ��������J�G���戀�N�q:�V�;w�j<N*G������[q�Nj�s��?�[���)�yg�@���@��S�9��^�VC�E�K�Pv
��6?�Z��Z��+c�<DU-w��?���S`�MdJO��8kj��5���℃='V�A�[�������!19��W|�[:X�P\��+����4�C���#(�k�l�[܂��vD����4�#�R9#��&F�fR��%�kj����r�����"��E�B�gꔀy�넬�w��k��� #C��c1����*,�M�(�զ53@F���nϗ).����+����{��`��ӡdc%|ަRz��9�/�XoO$�vhn�����J1�ޏ��p8�ӿ��W��R&FK�l�W�zt��$A�4�"���?�Z��Pa�\?�-y!u�U�o#C�KH�л䁔%�]߈ў|������J��E��p��Qn�)4s�]�u�0 �5����p3�|�:tA�Y= �S�3]���qo����<Ԅ�/��H�׎�߃W���^�7�Om�w�{����?�-�o��r����ف���;�aZ���	�@������5.Ǩ��w��#�u��;��K�/�Y��t��ne�Dv��"�:�$GX��MI�>F���ɰ���HU�B+���ݸt*����]�6�%o�HvrUB|6YB��f��ú]Y��r~ނဘEp�+=	eдO�����1�4�c���T��r�ҀYp�C8�!J�%.�l�U���cy�3��F�>jih�!�c�o�����@�?-��O\\�;X��η-r;�;�l�a\2���}�fA/J��bU�苏�G�M�3b~�F��f���ǹ;s�J��M�.��w��8Cd��ʈ���)3�&���C~���h+��9M� <��2D��ӣ���j�S��(�9a]�L9jXjj�V-3����ډ������_�յ	u@&	8��bM��zߐ}�Z����gb9 ���>l�yr�e�KjR��+y��m�>
7�����?�َ�:a�� �ESG�� ڭ�lL
A�Fk�$_�h�x�B1���j2ѿ��4��`:��9����0(<Lo��[�	�}��k��AY摽�3�E���6Lyͨ�z�+0�E���� �\�a�U�ѫa4s���khՕE�'T�8��s�]��������!�)s޲7�o�]���z�Si�"���
u�y��	�$�-m���� (�� Ex�� ���:�P����tD0%O.x��)��!_�Wd�z^诣[z��'ٻ�ȓ�	v�J�����kO(3�B�w6����vC�o�m%!S�.���|T��[�A�E�L5Xk[�#Ϸ��fb0��ˇ�r�m�r�PN^P�%��xr���ʎCP�_���<�u��v��+d����������	�+�S���l�l��ׯ�UY�3o�B��:��,6똠���J�X�i���;��u�:g!9t|	� NɊ���{�C�t4�
��̕��/K���o�W4�vQ���Z���n��������`�YG�Ot�I���xH��eOn��0f�2Q�!���OD��P4���ǥ�����3~H2���ú�|jL5����.����8���Q�Eo��@�D�x4�������<�]Ԑs��3��`�c��w����;��v����,��'s�c
�h��~2�O�ؠ�S��#�F��mFF�S�R��?y��B>$���NNjP���ÌƖ��T�jR���q��Y-Ojg�&_J~X�wɫ�]:�V��������h�'�y�I�����ִ����'�o�Q[C\�A��whϋ=2j��6qro���q�pK��_�̙ň��J��wgR���D�4	�Ӯa��a7*{�`qm�K�)K�����~�!6���q"���i�k���*�Z�e�*3oo��;�K�t*��?q�>&�;_}6�6���vEd�9���u�[�״��6#��;�.~(�Ѷ���-���R�o!�mc�dp5�=�@/�˛�� ��p^<����2�]Ж�V��+�*��?�ǀ�??��K���N�?�IT8U��=_j����5�	:�l�������U�3J��pU�)O���0�..D��z_�O����vQ�bR�A4�:5�v������^���:;~��޿c�S���ҫ;i#�?�%zk�,9uK��h"�ny��m�Ь��i2Tz�"�Z��x~��s+�;@� �t��Ν�u�.���;���;���d�v-sD�K5�Չ'=�L�d���\�3t����L,���ѳ��P�{�Y4M'{��09�<~XiZ�}t �̭�-�����ju�@��v��������6a��Q�����)h��b��3fˏ��2�58nq��A�NA�������*�̺o������PS�PԎ�,j��������f��;4�T��nT������+U`�HT���Ci=
��mc���=����g�����"���6���»���>�8�l�q��a��� ��*�7��)��*edy�$�o��|Vl���kuEh喣�����i���>�d7����ѵ����fC�j�u�GR�VL��U��-����)@$���J��l�F�lf�Ȯ�\\p��ZO\��h ��x��	C�$��*�!^�o�
��nʋ�U�tΖ�!c���]AKK�mL�[��ڵa�<lQ��)�}��Rc�|#T��k{~xjk���s��i���~��Xưh�31ә�9��N��ku�#a������aiYi��Hc���ǗF$�#��#�m5E�mh7:�����FY)B���a&�KY:�7���?l[���&�Fث/��+6˕/Y#�W���7Q0<3!�tuGQd��%T%`)=[v�]4(,�Y�y�Zr��9��c���'���������5aS_i�A��egFj�=�a��y����Kk�;>W����Y�-r���d�T}�u,tT�o�v\�qfut��yw����Q|������}ǉ>� %�|�\ {�2w�
)�C�)�L��,3�"$L`�Pe��	U���������('y��.��tdm�al |�K�ɋ����<U��j������9{��3��� c�����P'T��9��Z���u:U>}N�p��K���#���u�'�>aF_b�2(��\3*�N��5��z����,�*@+�?��C�X17ew���l����5��8���y'�(?�E�O���{�t��:���O�Bq�__����%u�׽�E ��^��0C����k��6��})���W�E+̜�f�7�2�C���ǘ��&Ked�u�So�&��%��j3m�JJ>��a�ms���W��L
��8jR�N�����>���7��u�S\��m��� �.�d6�oB����&W�>�s?CL$d�.�EƇ�)�~�!G! ��ݵ��͘%E��f��]7�z
�{%����=e95}��R��u�H��Z�s6,u�7*�|�<�"
lP�3s�C����#�1�^�`�a�4��=.½�eՎ	:�c����i3�n�&��ۄ�x�1Z%]
�ž4$%tȖ9ER���,?��T��ѳ:}�6�s����R#l,����vj��tZ�D�k�e�a�}�T���!hc��0��J��	^���/j����4��FjH����3K�i�*�mH��ҚcCwj��:�3r�˜!Q��M��>���v��fb�v�-o�l��Y2�\�,�<W��e�Ѭ6[s��V˩�11�4t�$��K���EL&P�*V*�?e�F����Gq;}L G'�mE\ʗ�u0�v�_��zA�ݒ~<�X�(>�x��w,�������Z�p�N���_�C�8L˚ES%A�w�j6�f���1�	{p���r4H�;��En����|��<�R�����*�����a4�ǅ����ɃV92I�p�=1L.��k�� ����'��P,*Z��m�Lt������-�A7�'��-ƒٶ6b�����<�����ٯR��x/�w*@re�7��3-�m���]%#_o�9q�k�C���j�3ý��Ɔc�)�Ŷ�G�O�ξ�����y�,i�{���}�u�/x"߁����F${�h/L���������?/�(�P�� 3�ۻuR�ոG���v�˪y��o�`���h���Kq��[�D+�;j^��4;r���D�@;N'Ge)(H�ˁb�0��y�B���r� ���t���m�O��*��?ܶ{E��a4U���V�Z�FI��z�U���m��rw�(|ܷX�rl�e�c���v��vZ1le���u�B��)�F���2�$*�d�L��Tc��YҊo�f���SW����A�Rh����++������(t���A��5�j	o�ba��-'6�Đ"��S����s�����U�-%��W �D�>�fG�`��]�BN�eC{���v�=g�B�^���B� �S�Σ+�/�J�s�|)���cD�	C�����9���a�G��]������O���U�A��ɏ�{+gMc1��U9��|�����߯�~4=$q��=���ȋa���<Qٝg�5��U��a�;�B~�7#b�Ҍ���tМ��
�T�Ӡ��h�LYPa�x@*o�D�5_������M�����j)�:up�L�o�x�=1ʑ5��zS�A>�^t���;K	�a7��C������K�y��sm0��K� {�9 )�{��������Sbt��~�j�v��54��������Yȡ�n�pw|l�U��{���2h���lw�o�&+��g��z�d@@����Q���㦩E^;�G<����q�ӿϓ~``���پ�F���ڗ6�W+U�
;wVΏ��P-�}1S�XU?�#��2<Q���
O���-�/얺ڣ�+��m�5�BF-���[C���E��U�US[#��W;�h��	��y��m�
�,���ڕWH�Kx~�}X���eE�K���/��JeFP��~ZZn/���;Ƿ�@vUY�/U�,T��d.ՠ6�0�~C��P��ѿ��`�"�L~��Mt��if)877W�v�������	s������GԂ��pfE���À9���c�ӟ��W)��\��j�(���{:�x�
�skƖ%�5�R��p��n��q��F��\/��o�3��I�+6�n/>��� UB+�׶�l"�{�w%�>�3���:jj3+����
��Y0�u���Q=)Y��ɔ��|�v��K���ӥ+ݬ���I棫�g/���������x��˯[#�#���F�'&<��K�yo��߄�{Q;�1� ���D2�H�v����l��Wo������[c@�w�o:�_���dr+a8�{D���5�j�����'6��� ���ax,�k%�6cX���9919�A;A�7���'��:���59�ɽ)��a�3gvl�Psu�=X���HvbY�e݁L���_��/v�Ƹ���>��m?��)���{��t�c�
���?��Ark�__�S���1��V�>io�E۷w��H��T<�v�/o��`�G ��t �M;��kp2C�Ҕ�`'q�hɞV��B�,��Y>�l���bHX����f�����t����S�m�ʒ�z�S�����4��_��g�ߺ�������~�(̅s����%�g/� �D�N߅�{����mY�N�t��� ʡ$y�������v�����@�эl�{�6��xW�ijmm�]厐�ŋ�����ɏO S�/xM��@�̮������A`kkɰ���$��9��HK�C���f8fl�r�<�͆jy�=X�l;�y��w6Z�a���f-���9�j]�_�t��ܗ�K�['���̨��Lq�|e�R�I|X7���B���T?:��"܅�î��S8��~���w��%�u����YК\Y��m-\��	(<ˢ�_J�>��n��Cy�*��0ӡ�X~�V+= �G"����ɿ�����@x�0e�I�������i����q�k^�%S��z~�=�j� �}�%���t������_l��p�sr�P.����;4�0WȒ �_�r��[?Rc���V��Wdx�=]�J�8���9��b�<Ֆ�|���s�2�pߋ|���r�nޯ�l߉�+q-��&��G�X���B|���>0�fZV�ٌR��ӿ��ph0��F�����&�$C����1��L;k�alr^ME�Wq�H�f {a��Ҕ?��WA��Cҝe�Nܹ�x�ge�o�7��~>�����g��6����k,2�]�"e�{�{!=�#̝��q?B� �*܍��L)��`^��"I���Dԟ�����]߾��Ҭmn�
��E��Er;^�Y|�N���+�x�V�<&������ں�
���ν�R&&&Ie�	�o~}�`n�;������N�s:�x��.���b�\},E���얥�����?<1#{����?�h���:�L��K�N����_GG*�����M!���R%d��Y�ڃW���؄e�$f�����;'��bF�^�W�V���$��ꯇ�[���:e�:4��hm����L��[���}C�l.cZ!���5��[F5�e�Z����\��'��nמJ  �x��R��VRE�ČcG�׺]^���y:2�h�`C����>n*LB�j�N^�e;P�Žg��gM�A�xP�I���Vcn��/߽i:�.�P.��`�.0��3{�5ɋ�ݫ077q�c��{/�T7�����:C��xS��J^��J��Ҽ�/�pN��u���[[�4�Т̫;i����D\�4vj�.�5��qF����~X�������ގ:��fh����3�B��x�?�;]8{W.�������<����ޑ�F>%�h̓F�U\RO����;7/-����jB���sF;C�P�~4�2�����ϐ`��	4B�ܸ�&�����4�N(_���`��yo�P�^D�CQ���6��"���=��rT�c\��k��Q?K�{@S�F_�Cg?L?�Lu��'h#���z�����P9�- ��]�ޗ�$g�{l���Z�����6�(N�3�9 );wIjW? p*Y�{�*J��|iQ���<���У�U����i2�%d0����0���?�����;��	?��79|{�cb����\� �����G�#�c�E�u��:�g���V�b#�KȪy�r�E7x���nW$[ ��i�O��������R�C�_�T��g��ɺ�~�v�� M�[��g^��3�dJ́���@?ϡ%6@c���@����rr�ޘZ��;�?;F�����҇Ǐ��ϝ�|��?����l�d�5f �����..)qb����(��[b�$��͖� 'i���E��p���񙇞��t
���0�������R����k_���}�����JwwzI	i�.G@@�1 �A�C��nP�kh��wo)(|���^k��x���&���݃���hw�W��j����"=�%M�"�|v��M4)Z�k�	oc��?~$����ct������a�D--XH$gDR�$3�Y��w���ޗg$�b�}�g<�R�-
ߘ�������:^�Uh�������2Rߧ�|扦���	ڰ́��{_rd���'��bœq_�8:�.C"��~F�����r��QP�0��f!�Ԙ����h���=[t���[���=@�������b������@��\A�Sg��P�6��I�
8
�	2"�:R������
�^���M�R��~n�ۛ�(ݕhF읿>�qC�k����blZ�3�?$^�"�V�X�l�kH��A�l=��&�6[4=c�_�ܧA�jy-o��X&�]��9�5��('#R�NΧ���1�
�;�q�;eX5�&߬s����B�����u��T�L�ݠ0Æ��^�⮶�}&c���|�;r���wx���xd?��P�J�1�]��:������Jb���U_1q�D|��q~`��c��=�"��kK���7�������8�}�*[T�e:�3Ͼև��+ }��Q;*���w�e�F�Q��x.P�㔢��ã�����®�P���6X��	}�"������-K������
�����K$�WoA�U��_n0{+㡳�����z�ڽ�"�A%[3"�W$I½��N���JJ=�/M�Xs�Բ�ڍd߀;�y%�,�&�2���	�%GV������+v�dڠ�̲ʧz�����A�9��:�Ѐ���$z|es�)��ƹ�����K�z�<�6�I\�qH�������*:dk��t��M�"SF�_+v}�E���L;C��R���
'���9+��qϡ��HIƶ}<��/^�bt�445��p:NR��`3��P�������h0��DAS�%�ѱ�W�_*���RK(s��f��������I�Z��f�ծ�����58�I/�����e
a?dr+	�(���X�c����u��L�\�,���ϖ6�2?]d�A���C��垹:"�$�}o���`��J��B_�X4�z�r%�F�7�}�_=�!>xtR�w�S�R,6���!;e�Ca�K��^����P��볅�`��?�z�⢰:?,�Y�);��:�eE�V���X��8m�
H�f�J�i�e�M��ÅD������6���K/�j������+cdX��]���ӝ��R&+�*�h�K���j��(���om2�)�r�{�}���'�wj*X=:-��������0s�r����i�Y8')�X��W�@�cp��U:V(�0����ՙvF���T1i��%I����̂�F�U��	5S�d C_�w��t;xI�e�v��y������]5��.�7�t-�:�"�)C���H���wX�W@Đ���7 9�VqI���QE���8.�=���9��ۀ�{���*&��T����/(=4��g,� 5Y
��V����NY���<ǃ��� "Bٮ�`�]余�)�?N��O�|���cl�Z����`�nZ�Nv���$���-�5�qOYJ(���`-����>W 0������ܓ���>@ͣ���Gzm2(j�
�,��R�e�%�J&�?�q�c�}���@-��h��p�[Vl��.qg��hΑ-���6�S'�������B�w�z �3�6c�0wr����Lkg�7�Ռ��!�nٔ���Edm\@��!���5�L(ڏH�����c��A�C�%Pp�(D�+�Dh�H��#�y��zb�ٙ�+��D����B��w0��Y}f�Ԣ���pˑZr�=R�P r�Ғ񂓑�<'OK�lD2̮U���к/�DY�DaU9����O�u�t���� �v�����;Ipp�[�I!����ZH�N�f��b��@�������5���>����+�aI�窫P+��M�X� ���Ǖ]BB�]Y���iՍ�&�b�f��᥾^�����Ó����|�bw��썇"B�r`���(�4M��&OdOE��Я�D��@p!`����:bP�Uf�xc�?q��rMII15���r�;�J���4���Q�)'	.]���7�D�d�wZ	2���=ꭷ�'��K3^e�Q}r��e��;��E���M����+#�<̭����n�R�r�ƈ��$~ZY��h�~�q]{��d��О��{��{aߩ�>��G�lv�]��U�iv)�����{�m���=)����$	 vvvT�*du�\٩����+n� 6�@�"��2j썅����Lσ֙��`4�W�x!S}��+�6C<��,>�v"%�30%�����-=(E�T� {�8nV���e���tG92@����
��ʈ�_�M�`Yڛ���J�"{zx���^���w�{�@ʿa<��Kj��� ;�k�ϼC8�R��,�:bd��^�>���Y��&F��C�z���N�Wb2��e���.���q����N'�\0p.@���E%|����E4(L	��E��<����h�ȴ���̔ߘ�t(�!Y�F6�%S=E��G��<�D3�8�@���k�T�G9���f�m���Z�&~Gq����@!0�{DjV}9����D5���>�8|>[{��p����o	@b����(/5���etר`j����y�̀
'�cT)~�y�6�����\����U]��CƝJJJ���$ѹ���ȯL�<��tX|�]��-੕�v�ߎfe1id]�V�=����Q�*�S�����|@}8���G����R���hh<����G�x��+�F�Ӷ%h�]7���ςk�[�?�K�����f@�����	��i�,#�(=�`�n���/��,��>s8�%|�-fP��!�z�H&���4�4��ܷT? ������G�B��oqZ=�'�:�k�OrQ�SE�n�x3z��!�r&�5���Aa�xM���s�/	L`�M�J�+/,U7�b�� Ѐ@L;}��mΣ��!��Yڝ��
mh��
����!e�^��0��HMM}_PP��� ͩ�1b744|w?�HQV$Jdiusp���ә��2�n`�X{@�6�7���Tт'n;~����c�� �c���ci~�o�d�7��D��tMi�l��|Se�7��]���͹��{�RK�(����L^�n��-ZZZ�**�6�oH��2H��nM�48^z�7����xL'��0E��GI��蓘����HJ���M��\~��{�� �d:،f����)�S~��M�կ�Y�nX⟄)�W�nrss{��jy��Uz�n�E���(6z_V$���{�9r���� �wn~$�)����>�=R�=���-�q���~5�S�A#����^���~���8 �vG�NN\���+�^y���e)$��p�`�����=ky�o����zz��W-(�1kCҲ߲�,�V%5p!φ�%���mE���я)پ	(��xt4ߠ��l�t@A�����BOjyO���Ȗ�`��m!��{��!"_@��R�~]�=�yߢ�?*�HƘ2������5���
�ˉ������Ὧ����P��u���I�&�M+}/V��(}(�@wV���݀e����z̏�TleO����iH�[�2���i�b<Kh�vm�C �S�=�,��ˀ�х���D�E��_S��:� �X�CHytYJKr���d��P�S1Eyu�;��Ç��W�m��64{�ۘ-P���*[ZZ���ƛ�`o{�R����«E�#��3+}k�W���,�Tm�}]H�8�Iż�{���92/����7莽opP��Lr�~���!�[���פ(3�ST�a))o��N���5WW��`��z:ӂ	��Vh	�.�@xWŲ�4����/?"�Xhom	�����R��*�KL�-�6�E/�%}�O�Ԇ�*hj�T��@���g�2kRU�J�_z\OC��.$RRB��]v����#���H>c��)mn��9�)�o�TJ��z�-�B��c�֋��a{mٟ �=U�t��o���Q302�}	ֱ2�{g@�M��^"���p�Q�a��:�}�ԇY�ލ.�1�a�A��<6(Fx����Z'�\��"�g�����u|ևi��J��/~G�9�Z���J�f�qӚ��?^��.���t�?�S����a�~_0�f��P\A	@}���Fr�Z��ֽ��vWZ�M�P4�Z6�16�b��)��Tj�(I�g��<s.����%m9�^*�V@�ϑ��C(R��Zi���.�����Tg��ER� V��_n㯭�9�&�	jT"%�=�_>�z;��	�@��"h��0�����Y����C):��P����3����F~qp�T����?�T��U�����茚ø�W��P���L-��W���y��r���fn�ڣMͱ�:��Kk9��0m����ʯg��l�����+D��[�鵻�ĭ��7 ���ߡ��e�'�P��|�r�]i��D�������o"v��Tg�yv S�~.u�s���Њ�H@����
Q��Prb]S�n�����Wy��ȵ���?����d�J�z�+E0,�����Ç��O'���̇g85TjOeM6�g�T�n}[����E�R�k���c$���ec�G�+
ëd��|���*tԲH]AX~�=!��}+'وPʱE{1�؏�/���ϣ��e�Ԋ�h�I�
�l�U5E�s_�<"h� ;hnMe辇�E;��ѭT�5I��ϴЭG�ٙ~��>x}�	�#t}�өŭ�*4���k�Xw.��;>���
/�p��_*�n�7��]�Q��N~����|(���PA(&Q����w|1�n���㨏���gz�Rq��
�
��l4�:Û�7�eF��E�ɐ���7�;���G�}����TѠ��e����x	���p���#K��	��r&���-|C$i����<�t��O n" "��1����@1�����
�c>올}���Ľ���:	ɝC��I�5���@GET6wҺ��9r�XǮmJ�꣌��˗�{�f�Ƶxo��#�����*�������Yk���R�����U5q��R�
/�Ө%##�`����`�z\���݂EKZ�O6D�lu!L�M��V$����x�CT֠�����6V6��������$���s��у�	�������a�k�O��r�ѴyBo4X���>���!���7���[H���m��~����k�ߓF�-
R� ���ǶAE��T��?9�ؐ[�z�w����̘]<<������X���_?���T�.���-nn :��i&H��&�xkS�"dq=����B�^0�5�	iP����1�o��>�����k�]]��ͅ�m�{X�Z�+'<�R��GZN
����ށA��om����OL�*{�;&؃�ԙ�������Ap����rA"s"9c:a<{Q�}_�쬕�0�~ҫ�0�(�8F��~q����� #�I�!�����e꥜>V��~8�b/	of)�á\�|�~��䉾}<�>�Ӭ�� ��v���ɁK����J8��O�NMͻk G��#��tG����#KO`��
��Q���by��p��Ԓ���uE��a?=Ռ�b�{O%~�[Zǟ��
�`_6_��#�̣4�HuB�v��:�-�����+|��+�~��������o��/7=���:<P���)��Ii��Pǭ������6��?lD�w��w�A�Wrk'. �NLa��Dm����թ�K|�}���2�F���4p�mK[b������K�:M��(� :���"9����F��7�Y���7��)�����Z��7�ޔ$?�#�����f�����e)��2�3��Z�y�Q��1����ޅ�����[���?���u�p�5-S 3#}'_�M���8?���waa�ws�V�KMv����b23[[�蒌nh]�x��,�O��;�RN2�-�N7'�VB
�
6w[E����5��/'�nb�c����4c����Z�V�j��~�6hƤ6!��N˿b� �&�[0���PNQ\{!��c���6�v�ފ���5Ķ����3��x�AAAAgxRy\%Jō��v�������Z�SVG"�
7,��"��E��C��Uￓ`�� ��7ʾ�l;P#J溽�r��_;��o���]�W76��˨��;���}J�Ԏ�J�Ԏ2X�(:���Sό"��'���& �/L �l�=t��6rsε�$Eh��Uƺ?{�����7�Ox�Lf��g��F5�ǣ��l2�Q������| � (��)���Oc�џp����p��R!��|����9�U��ڵɚ)��i��/Sx�s�R�g�M>��\h�Kw`��8�i4�˹U�A�u����sҊƻя�Ǘ��A�����K���s�7$�=Gw�Z�8��W�Ο��+]�k�$#"���x�	��3kδ
�-\�5A�ta�3o�v���`�������9���Qy�cN�tx��n��>�	@���N�
v1�l_"D�B���x�|4��V>n�Ί!E�y�Ԝ���kLfM��/���K��C�ԧ�f�:f���"I�5���!��B��x�Nþ3Ê{A&r��C���:W�[kICEy ���S)Gw�Wܨ�����#�U�I�7���G�9F،�G��T;���4��}���좛�8��&��Azd��H5L���TNR����g��������E�XQ��V�I}��B����:�r�%�Y��A����ӷ��*�x|�K�l#N#W��1��t}E�¦-b�в�k��O��;�Z�����!^�`�?]Tm�$�DP�z5xS���RX�ey_����˅�-屪�,��4�(�Q��_��ZBl!(�9͎���;�OLq�K� �~�� ��S��mP�<4l��h��Ol���O�A���Y+�x����/��(���^i�.�> %��և��4���L�	�EtRA����X<\mX�I0I�(��7��o�+g�
��|oS��җ͏���H0/�Ν
G�b?�8�����HA��O1�g������x�y��'W��"ܵ�Xh�U�UQ)�2JMo��(3�ww#vv�cx�f	��Z��,�,-��Lf�	���RYZD�w���Z�Fg7������d�N�j:��0=z�����
g7��g7r������eH���DS(��5l�E���U�)����e�q������K���9Г�}~�����Y5�Bo6%��X��Ǘ C>��|�(�̱���TUEz:S�Y`$*V�(�X��z_� bW�K��\Zw}�/;٨�V6������e]%Ӳ�x��l.�����)<��І������<�6�=�>�z��笉�W��X�Պ:ch��ꑽ�횝���b;,��5����F��L�a�&"�Vz��q2��6�y�]zn~^���N貕�t��h�"h1�<��W�����`m"�]M�/����R!x�����'�U'�/^�H����}�'��~�,���N����ѩ���w�/��D��9��a��<��K���hS�i_v4���� s3���(腘��6��5��9�/��Ld3��t����a��a��l�s,�\`���%������%~�����TUU�g5F<��{�}Hi���+�@F՚�W=	Y}����%(�F%�$�F���ߗ�����^`}�{�����|̚Ǽj�(�XWn2m߰�0��5�.�.��u�U�w&��෴OߜV�`�tʻ'�e�S���Ҝ��q9=�cQ)��C�q��v���$�~(�K�q�kg�>|90s<ALF?�m�NR䚬��?�"�(��B���&��ƨ�o6[��G�P0,�e�6�tEzߴ�&@~ޙM�|s�=�D��h���Y���^�t8�b��ab��l�2��ţ��c�E����4򺎉&M8;C�.�E��D6^�������n�� �G?"v^���.+Ba�QZ�>�,� �W�Mv�����:��P�7�׉�3��漌.��ݽ�1a3>���}������{�d������S���r���=6A�3i��f��~Ղ��P����`m��1|{o�x��'+ʮ{�[>�4�3\*��-���i'&� ��*�z�<&Z�K�t�B;OK�x�4��m�U++{�J$�W[`�8�c�(h��$Ƚ+������Y�217o��YM���D�z	��M�*�r���ėo{ʦ�'� ѻ㴎�&(�����!��W�!ɳ=e�ؓ?q�b=�(���2j�A`������(��$���S�Ο:;�ǁ�6&�e �J�%�j#�`(c{�!Q��y���<l��p&S��h�&�oڋ?؋=�ON��y����csll��o�S��Y=��w���rc'�7�7Q�W����㒙S��W��K�L����`c���~"��l����6]�e������S���;���_��s>��O5����<e����?�׷J�W�5��
U#�g�˵�kꪵ_�K�[˄]>/��n~���)�]� ����W��F*]�L�aB�F o��>Ժ*�T��X��`��礊;Jleee/g1����-Ѯ.����Y@JW|HS]]]���a؅[fm䌒�N���aՆ7��U�1S$����]�Դ�$�v%� ��ǇsK�T>f�^�s��KRB��������R����=%� :��?���]�{bӘ�!z�n�=~% <U*)ruu��l=\��@ik�Q{h�&������1�4_����
� �cm_��g\L��T��8�lो)))�̦�O�t�m"���+.T��7��ir\+:��1X;�&�Q1�������q� ?��8���������ŷ����\~פ�!�Rk��3l�5��F����#��)��*���@��qeĬqkD�I~"���![+���
2���y�y��#��;�Z��O,,,���Q�u�S�!���S��'	&�}]�-��%o�����h�E!���q���lD:�*�l�?.]-h�Ф�!�IM]޽���v0��AA?�n�w�;]O�"u�&۟{hP�w�v,�6Ďj�̝���0�������O�=s��p���˗@�״�u�t�Lک����ħ�W�=|||P�?�ݰ2��Z���e"+���R3�x?���i"$9<�<�U�b�'�<�9�J3����Uݨ��S�dV�G�@U58��0�M�ՅD֎"<i�����b�Ȉ��4�5Sy3�F���g�'&--ͤ�E�P��|�eK��9��_�2+�W�'%�����s}FJ-�&&&^��s{X��&]{�K�ǃ���m�3�_���f^��9�P�d���s�D"#AYm�U���V�>G��Z��j�<�W��_���|1v���,���I�m9PpF{܏ZZa����o�?ȩ��gM(.;sP��0�������x�� \�y1��]��~��I��{j���Κ��2���K`�m��G����nZIi�s?W���(���z|KTA�\���=_���`�:		Iv�>�?��KN����\�ץ)�*jh�3+���ȥ����_~�i��8�s�{��f��~R����+�^�Q�l����Nڶ�!R�B�f'�����&wyy�u��J�4��4«3P�����Q�V���ӫ�����~��Q�N?xk�Vض']=�ai49%����o.��ݭ�-A*z��Z ��<�%R����Q@0Npm��_��?,x��.S�����(@EEXwӭ��츌�g�7�T�l���ƥ�Q��=�0EԄP�o	\O����b�(`r���_f���#a���R	�������GTx����.�nk��=^{��n���GY���sq������I?:�����G���{����������{=�����M����'�j���>�6g����蹡�S�5���Cc��g�����'E�ޢ�������O:�Q�7�}�}y
z�����̇ޔx��
�i�6�y��Z۠Uxf�*6bp��t4L֗f���ϢDGC�:!X��Pl^(:J ���#���/�ټlhh���h�|��o�0�.�Xc}}]�.�e
~��g��t8�����R���H\�R����;��t0���`��@�4#�PUE�xZ��y(3pU��nC"	###�]�����XT�Wk���G��Ơ�k��Dhbס��D{[[��d�dɍp^���R&B�u�K�q�]x�#"3ي�O��$|=�j0?�~i�2���+����kX�XSK!/�`�˜�m�s�}\	�>���p����[1Ź's���4�~������E�f�V�	\�t?E����>ań�g
@sىxL_�����{�� n(�Е�T�CQ�W���	���&U����S��uR?ʆ���~�����.�
��sU�������2��r$�e��P2L�V��?�$�:�B��;�S�Oļ�HŢ#<թ����r�r��[he���LH�G���#6&H쪂��5i��^����&#��9>����h�$�*������T�1�&rb4�x"�}	2�sQZ7F�B�S�7Ot������x��i�_~��A�[��Cl�L�k�*A����ԏ�~�(���V�?xz�P�ut\s#wqh�Ќ�j&�<��	��l�J
x&���V�p����T2��+���BqS��S�{�_��&a?p/��P�Ǟ�<L���$$�O�P��J\���@�C��&
׫Ȁ���x��v�ފ���;��c�8��U�⧆T��֐�����I�B����� �F��,h,h����8j�`�ۧ�4��>�nʌ�y
�.����`���f�a��
�
�X��c�勔n>���ܤ]��s��e�iw5�[���<�>��5h�$�̘�ܗ�E'�=�ocx�Ƥ�2������P�`<i
�hb�}�E�_0=�E����t �X�J����+������>_��3'�l8�u���o���u��<-]<�h\,313k����d9��-CA����g�����gʋ����:�����l�t�\�?��h��^�;7����_Z:�����0
]��/}�A�7�ũ?V���8���LĬA ��ly/�QR����*�'�o�|�{FO��� P��8��t4i��������/.���[���i���H�u�5j�T������(��z�(�sz�������iQ �(��Of�~x�Y�G�⨮��������GmZ���-hi	�,aRfA+כZGF�{:E3�i��$J�c��w����-���M��X��n������~%�r�N��1�Ewd��p���V�~�{���|�gsxN^�_��v~���w��:g�<I�����P�^PSk��d�MK����^�i5H�W��;N��iwe,46
�`g,��	sF��9�R�m�Q��Q��QOV��ե���a---��g���&�x�b�7�p��WII�Z�I�kO����D�����땆�!�R=A�h���D��� ���q99�	����C�/��#㛂�}W�D�����o����7���{��VU=���i�����I���26H����K(v��Ҿ��R�!��us�t�y޶�-�N�6���޲�<��3wq�v�rm�?<�3⒚���
5���)Z3-�<}/a�-UlR r#�7o�g0��U�c�PSss��'2��)����Ϟ�]��@'u]�~����SJ��}W�����92�LƩx34>��D���\�UqqqLӛ)�(0�,m�����cakpJ�G}6��N��tA�P��ȖX�?��]���M�853���-��NT5��1F�i���f��<Ơy����z#�W�C�ѻ���O�����y���f�gk���� Dj
�M�ZRv..�m,D�\J�����8@в��E��\A�c��SI�W;����&�NFCC���asiii\n.�_mp�%���d_l��و9�=
�� ��85�c��?�eê�B���Ka5���>�.�s��8�����6&�W9g���pe��2)Ϻ��<I��܁loo�[緙�4K,�A�'Ep,�KI� �hǩ�����+7����G����d.͟��5��O�v�P�P�0m���5�B��""����i2�����(�J�TɉsѼ�ȳ)(S����;�8�mn��@��(�wC&%-\nnnjZ���zj�C@�(���.�~����p>���6Z�b����Y������iKKK�{�������׽��o*���'�] =��0�]�ob��6<0 �r�Cn�),,�@U���3�1N��R1��6�8��0��1(������6���\RHS��N4��%P*�,�h�e@��3I{Ս���V�X�b���#�^z��K������n�ز�J=^'IX_��RN-����S��3j8����k��iɧ%	6o�h�؀�i�?�F��\&&8�	.�F���q-7�ԣ��%��Wy��3r�Z4�8�/�#ȴ�ʳǴ�������Kk���T�( Q�QE>��A�|���Z�	Ý7�i-�[#�B�=��i����{Qig]��¿�:X�ߣ����O�_�VZ�k*V3+?S~���y��C{��1���N��`�T�H���3�[��������@���Lq._�|�{����Ւ{l�l�ݞ����:����~E-����N����6��a����޻/*W���9y쭣���~h�ࡩ;=�Ю��g��W���:�}��?�>��1�,��S�R�����(�FAR��R��m%s�M�����N����P�re��Ocxڿ	ц(�i\Lܸr����'��e�ɇ�>�stmj�/�^<1��2�>�B)�zZI�Ɩ�U����Q�0L}Z+�'LY`~B�$��wm[3O��I�a�f6f��ã?Ttu���/M�'�����Zș��'�p�g8���W.�i�+�y^=�b�D���~ׇ;�]+��5�і&?p�ZL��M� $YJ�x��ŋ��<.�>k�p��9QS���]����"�#;t�I�In�dE�bT/�q��h����"�,<,�=f��QB%��2�%%���*W-���K�dJ����)�@�4��[+�� �^�Mr+��_�����r!��	�S��9�L-�󮻸�� %=�?,:!H�GCrZz=�����r�bU���W�і����gB�Ǉm�T+�kt�1�X�7ì<0�s�����yk�R�M`V��MQ�2�a���*v��8�-�l w6Ĭm/�ޑ< _�h�
����-������{;J)�xG,���;�0����|���~�XR��2�]hh�5>����~	����%�wV�����<he�l
Žt�RnoR��q������˸&�����.���(�;���f�Kd|[���sۚ�6�&�Mȸ�:�]����#�����0�V�ɨ����G�sv�࢖=1������>{#pQf#Tq/J�Efsۀv��}.�8����\�L�C8-x���sl�n��u��3E�rN�B�Bk�Vf��v�>��vx%�R��/�ha.}���-M�i�,vA�i���G��p�\6=�|)+��3J1�MmT���𢶅$� %:��j�������C��2́�!��%0�z^#R�"�R���}�W��-����ԵP�yc(�q���8�����,6�;��}��R;���n{�6�LL�l_���PO����cY��D���&���Io�8�v�N+#;�Fc&� q����Z��0�ѷKwZ�[w\��ֺO)��ػ��D���Z�j�$M���4�7��Ё�Dk;L�U��v���sW/TL\ŒD��1��na��@��	�a�E^]�cf�����Ą��o��ZkX�h�<�tj�q(�雚Z�ѣzlb#����"s_6	��g�h⁻ʨ|,ԯ���>Y����¹@�	�x�no4�{)�-�:1s����ЍYA����g'՗��5F_<�:3&99���U�VA!�	�ѱ���{|B�w�gV�m��tn@�7�ù��6c����+7�w&���m���mxIC��+w�|������r�im>�@韭7���H�7
�?n^t��]JƄ𕃚�/��IJy||<�&�QM�з`=�l$�|�!�v�[���`ͮz��9��x�{�ill����u�(4�#�Zo��˃k��G�J��[�^-��R���α�J������3a�@�0d��~��_UKt��~e����W��b�w�5��[��l�uQ�猱dN��>{_����\��V����_I��t�pׁ����1��tu��jR*w$Hz��|"��rɉ2�թ
c�&�>H$~f���3��J�暏l�U��z���_��Դ@%4����1nݵhJ��7�u\�]��!��vZKINvO��`����a�������A�jod��K�h���t�A;5qqȵ��/�� �Q��D��|P>b���YONr��5wM��a�3���2����5m�|�CK�v���I����>E�ѿd)0K#�����$��b�l�+�Ƴ�s�Ό�KmP�7�F�W4�S��#+��U�ۓ���b�_<ǁ�B�qˮL��ƍҦ�6g�D춓F)[I�5������j_��\7'�-L�,�˩z\{���(4L&d��F �N/u�7윢��](f�*�c��W�5]��;�l�O[�t��1Bh�R���m�da�^�\�� �������r���cն8��RJ�Ȱ� =��\ ��^��Z���HM�������>�VG����ܖ�(RL(>�"��	K���b&���"w�љ/?�~{��.����S�;/G R��&�W{HG)D�	?bxtߪX#��z�l�2ޢ+�Uj�ϙ��1A ��gw`�="}�� !񽍁IZ7j�l�>�*D	g��	���ڱT�^IV�R(�W�H�b��:I�4�}�x�\���ꚍ�~�eϙ�L1�num5^F>������3��uɱ�2�޻��R�W	7�9�OZ ��yC�5|���w���`IC����XV����<���]���q*qM���Ę���p� 0$�?]S�����X�أ�(,E���]r���%�Q��r�%}T\$^]\��`$j�Ї�ߞh��!*�����!!��)|F��c>{�[��他8��*���0��/I>N�0Rb9�g��V���v`k���:V�VC:ʖi��B��%��>r�,�5�[�7i*Y�k)X"W���߳'<+�p;*�*�6�W� ���u -~�׆�RjP�;E�&�k6wU@�Ss��#��`ЮCc��;X-5����&�0BB��g�S��C{	������c��{%~�
S�!Y1Lh�!���
��fx�{CB�̰u��̵��[ޮ�,K2U$�����;�O���b��x����G��%k�8�������y�D�����.����gQ��S����3be<N���uxt0��Y��&�Zc�j&�vC?ڙ͆a�@���p��|�����`?�+�0o�``�a糀;�,�⊢�sd�W��F�5�@�%+�=���.G�S՚vO��X��˫5:���у���X�����#�+�S��L��B_ɗޒ;�gn���ڀ��a�`�!��iږ��L)�=����ޡ��TN-j��5{;�C��k���ǸB�C����3p�"�0�R�Ƽm�jձ�ݫ�}̽�ްf��Y9�N�.E��mX6�C�g#�]��7�݄|�bܟ��g���A�$��p�u=���@�W�.�,$,,,Y�[��i+2��G�~��I ���n�w�\��Zn %O���G�)-���$J����� 't���ٜ[q㙅|�پv�J��������,#����7����d��_�_�����+�U�k�P�Hi��^�T��i/���7{�.��G��L{��1�k����s0F�1P������L_�7�����c�l�(�!�Ѭ�/���A.����\f+��ॸ����l6@��!�l{K�1�?17w�?G"���@�O��|��	�S��,�-����͝9s&�ica.��t���w��F�J~}|+
�˧~��U_t=�k�6���@�$t�ڊ�D�`����}+Y�;1�D���e�+t��q��?�s�'��j�hk:��2\�l��z��^�%/ݶ��C�3����ZBU��]/�h��X��R�՞λ�ܿ(���nىbly��IrB�4bi=���b��ٜ��������1��a�{{�6�c�銱��j� �9[�2�HD�q��I�lg�bq]���"�>�1yG�]�����ֱ�!}�W͟�]�\p]�qe&�є�oJ�Ɨ6b~�{Y��L���"�bQh"r��@r�a �d:�%a��'FY�YEB5#�JK�?�7"���6�Uʅevf��Q��<gm}������Ɔ�#ȿ����;=\!�Aa�����9�9(��F�`�3;�\Cn���ηr �)�JY��
f{H��T�@���e�:Z��[ޟ��|���3�C� �I6fu�+C��w�t�E ����]@eK�
�[�@�e�<����cd7FYcع����*nXG
�f�M��
��؉L�kC\S�e��G3��>7�&-x�lXD�7�Q@#j�E�C���
J��j뮇����V�ܬڑ�����j��pp���;�A����ݼ']��Jn-;��A��E64�NR���.�������mv�ܦ��3M�tc����H�x�?o�QG���@�3q4ut
��$}��C��/������LlV�Ǎ����~����W�#��e)l�]�I�Y ���
�$���	���"<�`>%|��Q�P���66���5��P�H�Z-ƠR����ӹ<�����%-��r�>�4���}A*<��o�\�,����N:&M�	��䗓L�JR#���a�@��@�';Mv��ԭ�c"��j���PM��/Ta�;��ɺ��D.��jxɦg\i��+Q-���~��&´��@��T��q#�1].ɓ�&E�@�w!�$/D�Ƭ�Юs絘��d�ԇΥ����r�!/��ݽf���f,�d�/t7��y����O,���V��Qu��KJN��>=�;WWW]�F��t1~U��g_ݤk����ok�G"���n6���_��*�Z�$]�Zb&��ݶ[n迯�k�=6�|z�յ��Ȟ����_�R��P1v���y��.��e�p��-Ǆ�J[Su���S|Ձ�i�v���+�������e{rE�(
�M��wT7�&��R�b\+��MÆ�7�G�"u��L��M�$�����K�R88��s�D���";�F�D?���o�{�
�|���/�|X���
u��-���>OĵU>�}����� K�;���@(EM���7M�uԋ��=-N�����T~�
��9��:��`L-Z.-<���ɶ��j0��(~\4���|�h^�����v��!�jQTB���r����
�'�L}��{bpf�.i�j�X)^���	%�/��p��)�f5���o���L�Y2�	����<..��^���S�}��B�纳vMm���J�����ؿ�N�@�[=�2,���%5�߿T f�%i8տ��ޏ���!v7BŪ)�>W0�f+�P�!��$'���i葓>Oq�����
�q�i�e�����͝r�ُ}?���f�_p���#�r��v��, ��p�&,6�l\u@����9@B���!�!��-)-ݩ�4���	Hw(�1BZ��������W��?{�m��<�9�3�$ˁ�d��f�bS��2��99�Ǒ7V�Ő⠠ Ú�6�瓁�J��ώ+�B���Ty|�,����zAk<��`��Q?�ԶGgnz!�Ly��G�r�H�!�6� }��y���a/h$���鈛�Պу��]3�.��+��y��p��ן�Y�=�R��-�&�^��wE�R	�l����t�R��Br!����F�|� 1>�ߴ��:l���"���İH���cDvt�  $(Ȏ\q�k�{QM��olMl}�#�3_'<A���)���?xA���/_"=���������A�b��K�v]⩭�><�����o�^><q�\�M)���s����ދ,�<�)�Z	ۛ�������E�{��i,����Jd�Y�6^$W�@���l3�em�6��=�>R!�I�Pˍ��II-�==�͎ۨ��8}�RF�*�k��I�Gh\���2�R�E5�Q�E�r�L��:�<��3+߸�UZ�ha�+L�\��|��.G���0�&4H�4쩒����6�~��ģ���.p�2dddd�������n�W>�P=�V�1���=FG��=�G �,�<�^��fZ����zg����7������<L �z���˽n��ۨ{S�&`��� �\wW�	I��0q�h��dn��L�b�z�����&1�֪iXT����y ���ô)<� PmGT���Xq��j�9�Z�XIk�|;��:�WU9H:�b�uջ��"��U�Us]o��a��3o*��lޓ�v<�R�u����50F-�{B��*t��u�uxc?�2.��<���K��Z!|���W6��&�8[=�k�)7�|u�9'���)���m�)�!j��[��d�4���>B�N�%�z"�	5X��E��)�
D��i���ȃG��*�YTמ�Y��?�~&�́�hg�{��K[�_��$�10�^�*1l��%��e�"�("k�%T�x�b����RpRg=����do�|�)�\W~*Ӷ-+�����b<���/6	%01���(�^�2�9��[�~�(���DLv�`�^ {�������o-��5/�+��HH4�֙�ޫ����;�����Ω0�q�.Q��	�#o�-�ڀ
Hz	7͔i���z�s[�&ϫ;�O�����������5CÉ��Lpu��R��8nC�K�b���m̥��w7����xf03~�f	�S*Yϐ��E`�Ges����nr�@��.�Di����sԣ���R࿟=կ���i;J�Xv�E!d	�C�,�k
S�#e����$8��ҟ<���v�h����`u�#7��B����?�D �nZ��˗tO�3)WSk��*h�r��~~�`\�èm�+}l��?j�=����5p����ü�HP[I�������Ti���pFz���M/���w)0�6X��6�}����J^ޭך^����)-F��n�d�lY�gZ.��(�	,��Au�]-�i��V ��.��g���$�JmC�{s�c	jv�e��-{��狝��R����-oxQ�?��I�W�J�gֈ��h>�#�d�a5]{��h��Hq�WJ���=��Z*˵Ý����U�[�|	�p�U��q����dypB$_�lW�~�`w�y@�Ǌ��S�� 2� �H�����q�J��4�������Oǘ�C|� ������fr�&�_{��!��R�cK����N�wXEa��F&w��G��5<���(��pO[Q��)�Ә*��J#w?�t�!@��n��������-�Y�\ ͘�f��>e)�T�8�Z�L�.��p�����:�^I��N�kr�S���R"�;�D<<m|�O���]�Ƕ��򈛛��;�1�0���{d����^�*��o�N� ��Q�h�b��zg���<��,)-�xt���?�
�-��ߖ3���O���O��MV(�_f��&��{b2�چ>�]������|�^:@���Y��+�Ѩ��@ъI� ��$���=y�9��$��B�:�V;�a�S~�Vt��m���}OaAa�*s��uo�ρm:�c��Z�{Ϲ��vێ��6D����e�dLXC��;e����+F�扗�ǔS�7�'������n�^�\��)��@�=����UR0��<�X��e%��UU���*�BO�m�Z��N�g�~�z���eϢy�Jk)j��t\_�7��ͧFz����Q&т��\�U�e����BG�ߴ���%��˺�X��eR�4g�x��.�&H��(󣞩i�7�J`�.\f�S���ȇ �{����'����M�qѐT��'�[���ޒ�Kg9c4�!m�<��Z����B��Į>��	)����b���3�cnZp��>y��`,Z4���M^�ɺ���J���+ύ��
�hXj��l3�q�Ԯ��$$���b�{H�?�c֙��^R�]M�).+709,!��0�xy�C�+uۥ�_O<�&4�<b���;(�ap*�n�"�s!��^�Ek^�%�Cx���QS1D�z^3�OB�Ӈ.+�?-PiN"���?���X�v<���E�?S%%�_s��J�Gx|�,�@��}Ә��	�s��}LoqGU���������7�~��Q!7�Ã6�hݎG"�_�ݠ+ s���Rc;sI�<�n�3!��F�F���6J�3h���RQ��V�(K�A��X!Xx��ϧ�.k�J'6m����f>�EY,�8:��K7�r�F�w
�B,y�*�<BL묯�Á�%�^u������5�j��$��vf]<��.=��b���l�.��t��b��_�*s�sp�h]Jb r-��[�)A����U�����*�T&v��Jhn�o�e"��tU�cA�Q�N�g�*�ݜ�0U�9��WFs" |w���̶����a�bn�Yk9D\�@��e�\)!�p�tf�������5�[:P,(���37�f����`�GN'iդBGG��<�F�un�E!��f.ϓ0`�͏ȟۀU�gt�?�z��!x~��Vu�Y!��~@���<1�����MAǧ�l�:Ky�0˗ �9lO��67-�P8�G����n�S	�54������QM"��Y�]�sυ���z3�� ��U�����V�r��⦡�A�B�D4�߲�0�����IV_�9�*H��xW�B�l�d��i1���0zw�{,��+�0R��;�W�0��O���lm�
*1�B,~�K�|����-�l�TZt�i�W�i����R���t�[���FS�nՖ�q�xx;)͗���D\�tUl����Y��� ���œ ������DoT������Mk6�T�Avr��Bc��vŮ�1�'���.4T��m{뮇bi�u
��/��V�����>YS]�廊~bs��{�YF?B0��ER�ظ�����dB��pc��`��j�tenm�L	�H�_��m��323��𱕿�K�}��"0����WU*))�6�D{0��zII�PJ;�un��d�P&jj��7"�0��n�/��N	�U��|o��_�D�i���9q����n3��9L���CS�v���8
S�3}�<�*�kʐ�S��l��,�ŏ�!��w�����@Z�9r�v���V�8���>�n�T	8@���4���6hzD��¯��<7d�\g�Yj5�ӗ���k�'��RAZ\�i���(wr{�ӗ˨�iN�^��5X��,qr�:�Hy�4����㠭<��-+�O,�kz�XsJ�,�vz��SF	sUsH5�%==!��X�������1��D��|&������v���r�Pϯ��|4��Y^����kҷ�7�g��7���W5=��A?�e�vL �dYuzZZ�*/��ottb�����&]�D�ؿ�b��썴��r�q��7P��GS!�!e-���6	��+@�����{��0y�"�AX���k��v!`DEiTb^����Ez�3�g���Au������y�Ҁ�W*�ގ�z�/�_���@�kpC���+a޶��w��s��k-#�� ���
L|�H�������]ܸM��bo��d����
�O�h�t�I�b�;���\���{^�i��[�j�ey����)���
����au���,�(�A�y|\��j7'�u�C\��v��j8�--W�<LNX*VD���:\��(t�e{��jijR���1�1�"őa�q�k��[dPZ�W�%.yz��7`;O�ܼ0�������R��ٖ��b׻U�J�zYf�hau+L���EZ�J�0�#U3l���Bn�h1����.�r�R�:���O���Gݟ	�����A�t5A�8O.��І�8��6�^a��v�i��==�z���5�nx��@rNV��Cc�S��|:����^h)f�ot��.Xm���p�̅��F]���U���1�Vy�=b<�i]<1Y�R<Y�b�nk��X;j�мء����&��fM�E�%�=7e{3>}�����&����wb��Y�[���溦r�k���&o�'?����1C�s�	y�O2
�� bX�oO�9�b��׷��w�n����p�C��]�t-�u�s������(���%s�<{�g�R=�ݭ�*�Ճ�"�������-w�I��Z}�Z�tp�3�~�Ӛg�7b�>���r��K�J��%5�ո����8�K��,x�.n��6��Zp.�/�˓S�����Z��6s�A�-�?�_��U���j!�@�c-0&k�<�O"SZR6�Z0Oڡ��?.c���̛��2b�T��x��#��f�h�K���3M����E��a��R��yP��+����+����������\�8n�ê�r���+�����%�tj���~�����������٭���-Mi���%0�(�ђ�l�RE�HN��:���g
�O5�nH{���;��By�/����.�����,��e�wW��	ɬ'n���6֘�Vr���@�O��d���"R�:{e[z��S$��Lȴ�m����1�[cY9؍n>
�$�����>��[�$��s[7�w�{����,��i5�w1<`����v��.9JW\*Pd5<�f�D|@<{39ꐧ�i��� Z��hCX�O�M��fk9ű�|2������t��I������T��XŮ���P�B��	�J)7*fS��I��2g빥YEM,_�ֱ�*6m(}�s��g?s6���>��޴\9�K��:�:���c��g2]��"�:#d~�7�XYٻ7� 53�Ͳ��N��/X��>��!
xRo:8;i�Z�5V��w�J�}�o��b�b~���ɓ����.�3݌�")��=.��� f�m���/�a�w��*�Z��[��g*ىf� ��4���K��멫F4G�����O�v�O�X1�(�g�F��E��$j"��p����s�*��-kM�7F�V���J��\zW�\�d��6$�b�����>�(�MΩ�|�5n�ԧ��I��K��c�]��s�����0������?e\�h7�c�E*?�PE)�nji�����Y*U=����z����V?����pL���R��M�C.����M�ܧ����ΕP�i�T�us0A>Fm���c�6��.���11�[����w9����;�{F.����g�V���/)�%��.� ������WSݲR;w�)n�1�-�?b�����,hgiq�c�J�2k����X&������Xm3G�ʻ����{
�V�_�mV����#FS@p�h�=�����AD ��wj�ANyݸ�x+��ܲ�h���-KL3��n�M*�`޷ ��ﴢE0 ��V���zøX:�_n�R�#	�ݼ�6Q�%��a�O%��>��-��E���iEj��$ߒ��c�e�6�e�Qg4�5���d޳P�jܡj}��%�\m�A��.���9GGKy�-�qah�U�Opj;ͪ6�����E��2i�I���2V*��[3Z������I�轸�%
������ @�q�WfKT��V�Q	�����2�^��w<n���{*��-�v���_鎉r_)���\�ɟ�W���L�)�8�a�3�@��3Vn�ji�^^,Yr+e��' 6�/�4���n�;�w�8���3�#��b�Gm�3������u��#!��Xt�U����XQC ö"�,~��u���+Q��'o��{kOe�h�ŉ�������|D�L�)���!�b�>C���n\��8
��һ@��a�4y�q�kͶv�jV����X����L�aTk�C�L���.˾P��X������,k���B���}S���������
QTT��Z9%%r44G�7�WMt��Ϟ�;t��a|���h胸�N-}Z��޷}ު�)��/[u8���Gk�O��?��(+S�d.J�IZ�|y�-��q1^F�E/���Ϗ�oy��c��p������T���@��+o��{�>��{.%�y�'rT������}��>���H0� �ݫE��m�|��qV,
-�8�c~2�Q�XQL�Vz��.s���������.�V��n�W�{��M5�L��2'j�:U�"uD���rs�L{.�L8G��c�����u���K&3����YۺA�09�Z����������0ѓ�$��/��'�]���9<�V�Ew�DQ3NV�P���53��CU��ӳ
�ߜ��v��qnc���'��k�����Fl�+�#�\63���f�|��>畵2Ss)�d��2#���ʤB�Y���^<Ǽk����V��K���@⻛,�^Vk�H	�~�����K���,#|�`��5�o���>�Ғm{�B�4'�l#� ю����B8��� �pjk���r�<!x%9^�K�I�g�z6��#b��tQ"U����V�C.T��(]
�-'�ђ�I�Ut���H�YJdL����]���Jz,"m*���9hR�>���}�Y����c���T��0S��ဩv�OI��g����?v!�b|��*)��A�B��b8��S��[�N�����{��ՀF
���`���A�j%d ��l���'�̀Ϟ�Y��mB U9���0^�G��+g�����~�8��ü������d^�񓾻�&�#�r���&��L�ni��� ���藕E�[�6�WR^2���ϑ}����!��ָ)�\88�R���s'��gث�O[y.�c�M��f��X�%�Wj�/g��v�7[̷{���+�������Ëk�d`�	w@x[WAt�p�k���:)'/5i�0���iZ1_�*�i���b&�&���.�}4��;t:ي/ l��퉋Ǝ#ŝ��(� ��NkhQ�TϨV��D�J!��D��&!�����"fcS�2���ɩ�V���n�x_H�զf��-z���[���L�0T,[DT�`�$u4����!C�l�Om�(���9��^����k���
3�!bz���)=���<h�i�n-��q��uHK_�;�ƴ�_%F�y������4��j��u�.�7FA��iߎKXٯ3�T��0f��j�d^�oQ�@۞9����:U��Ė�����\*@���\����)Mv\�1���:��d���JJ��gu-�-��bZ���]]�<�Bc�0�ˌnU���7;�)��eo�a��A��J��}6�xSN-ejIF1HG+.�ŋ�긊���*
V$*`c�xz����1��s
���?v ��w0WG���]L���}��4loM�?�0�g��r�!°����ARz�AO��U����k�D*�����Bt3h�#�%�nU:�gB���'��,\�6��b]��~��JnvK!Y����p q�����O��	g�1�V�[?�G�qS�ZnOT��x~��2?����_Z�up�'��M#"w�:��PFH�$z����Y��w�a�b�]���U�F,�z�c<��!c�~t��q|U5�o���I���}��0@��"㪹�+N��w�k��2��$(��X�y��OW-Ō%Tq��������9���y�j,k�\=�a-�*�����`���7_�8>~a�g;7!��C�hÄ��N��	�����G�<zGN�:�f�.
>���< M]�W�署���,����ۧ�Z\��Ԉ�R5���''5�F�R�>v������I�����zU�e�$��Y����,��R���+1fRu������֤�/���d�)I��gn�$��#>�V���^��E�Gx&��M<4ST{��ߥ�
�Y�3W#�汝yG���c;4�p�"�&��aa,�H�k�U%���Zm�w��`�v%z.�}��^_�KR��o��	@B�
��`�����|�+��)flL�� Z�k�F0	�H�Q#��̣�99M�䷾����.!$$��<��]3?~��������cTB^��SS��m�g��-�\��2|�T�Ղئ�n�B?�kDœ�Ê���o���j��oج��� �
J}��γc�Z���{���QkNg��L�f���y�W�ߊ���'p���/�AroS��YHȎ8�PІ3��9��|i��oIr�(qHH�� ���2����J]��yL^H=�KO �Kk߄l���ۘ���V��~$�`F�ܥq�r��Og>�y�����������#4���=�ׇ�j��_�I=�`�]j&�k���b����~�G�+��p�Z�Q;Qy��J��{�~`t"իd�XfͿҩ7-������gB+�Y�O��?�# ��T�/����E�h�L����\�T`O��p��T��ڜ{�N0
p瞧��ޛ�������W�F����km-�m��z>�������!2g��k�[�6+�ۙ��u����?	4�}����m��CKT���B��'"xމ9���]=�M�G��y�ĥ�n��\=�3p��H�+~�g��ʍ��/��9@�K��+��C�#I�'���w�Ͻ%��XJ�"A)���O&<#6w�0X$ar�Mh{G��M���lY^q�9��)�a�M�#K�J���5++;�<`YcG��dq���V�~7��n�'��|r��b�����s�X���}����&)�Th�OW� !mU����eA������a3y�q3�r��GNmO��h��R�w�Q�G����ܨ�-����ՌE�fX��`�0\�C�7K���:D��8�1��a�ϑ���+����^=_Ǳ��f��3ՎT7��*g�p��{�F[,��75�I?[ޅ�s�"�@Ǥ��م����Lܜ8������oٮw;j$�)"Y�/��E���<(�x���%��u�_�Y�b@�����'���/�ضc��0��<��XUX�I�s>g���mOn��gWX�1v�42<ܙf��kL�@�����%$�HJH?77/�1$�l}���.���f����9�cQԶ�wq'H�� �����}��E����Y�Q�4A�x��?�H�щ��D��t!5��Gc�V�6↙Zi���$�iȑTy�	��u�{��XsYa(�įq�&���<���F8ڛ
_���M`1B���ƀ	`�*��j��*8>�+�" 1��ˆN�*'� m�t_�Kz�t��X�U�H�e�ԊB1���k�����%��[�53�|�6���v6����@ �7�r�m �	J��6�j����$Nc=Zԝ��Pޥ�!�b�������|is���.ڢ����Z�G��2`7H�Y�2�%0��H)���jN�eUh��
~Ft9�u�g�w �ӎ=�
� মS�p�Y�Ϧ�ڸ�ѣ��������S�E�te ���Y���5����.�:ʇo@��i�b;e�]�\j;z�q�q���͵��ˈ.���cF�Snn���<q��m���oM0��ν<x�y����]o\��
o�;p��햡�D�ex?���e��] ��v���EJ`��{��w9I���R## ���-=��80���
c̬F��&�p�m�'��(1�g���R^֠���*�F&x�e���NO'�kԶǋK7��.�`��1=�G�R�][�s�J����%|
$Y&�50�G���\XPY_���������q�qU^��/�$1`�^ތR���R��q��3[ �%��k�ߛ�~�Ȏ��Q����($eZ#q�JY�~�� ��!@�A6�]�J��p��2=%bJ���s�kѵYRw�ƛcF��12|Wk 6�8��.�s�Yo�iR>�
���7mhxPl�hADBc-��<�@I�wQ�J��y�Nq�t������q5����1��nx�C��\�nm�MC7��J��<�b��0���9EYII(,��_�F�@X�P�Vt;�2[�lh�a�E�̉[��~5��G���]8��1���Jj {�-E�^��]�Mj��A��&=�n�:P�6j��#��:7I����cl�g$�~����Q0$�^�NZ�撐P�2=M/�r쨡e��5����T1�d��a��6���h��-��Rk+%�Ch��$M#m=MN�vS*�������Y�]��%��!�ޠbJ������<Rݸ�����2�$��22��L���D �-�,��r�'?����y�a8{��*�P �A>���0��T�L좄8oa��	��N���AP�2x#*�ᶔZ2t
o�+�m@�|�Mд&C��_.t�౏���{�ȃ���(0nu��#����᧓�ҶV^m��>8���f��9i1(��P�@� ��a�װ,�gW�J��6�z9�?V��x��o���0�Y�bk��>�J�a�3ȫ-,���x*��8kĂ��ñ�����<���&�ɘ¬�~�&���*���
��Y�Q�cz����O>�w�냿o�mFD�����Eek~�|�$��p�)��)	��Z���]�Ղ����lM�.��B�n���W��+��N�Ę�~���9 i'ð��v�?x(Ml�l^�+�;�S�4QR�Rv�eV��P� ���06�WI�c�u/�-�^��V��fj
�fpoʫ�6���-9}Z�8,R��\z�������Z���o�S�}ԓ��>:�4g�g���\υ����� d/<�/�N�L�	H܆�������m�5M�ٔퟯu7�-�RZȝ�b��ŭZ v�8u�~��ƛ���������g͍! v��@�?��_���G�lf���=�2J�t��38Wf	�k���U���ފ�.@�v̖�qA�����J��'����u-������Έ��1���� 5���ܙU)D�收�0�8�#<���=8Q��8F��衙lx=?�ew9#��?Q����YO�;\]���j�l&eן��r����We�o=R_vQ�׆�+��W}ve1o�m��u}�f�V�N�q�^6%�U��0"l�2P����@�V�uœ�<Դ�/� Hg��нm]�5���[��gw�]a���k+f���C򾔼WBl �u���6��B]��Q����|�@ps߁&5��l1��_���\O�$��9��&Y��٩�|���T��H�@�`���T93�B4v��^���f�	ϗ�M9XETP��yCW
��6����2��)�y5��
!6��4{ {�3x��VLYĿ�TBSD6��P���=�F���ň���0Ȍ��;S��k���f$���F�%auo$�2/g�0_E�8X/ϭ���.��o���#8Tj�W��H�f�*^g|)�� ޝ	\"(
f�yrp8;��=JV��)�����7��{~�c=ZZ&V'n&_h����;̛������pD�,U^���ĉŭ�&ȫ�����j&=}�R�Ƃv��r�����$��K+�De��'m�ӫ�_��P1L�9�qwZ�e
9�<�k�n7��v<�n"�l^�+��#�A����/�i'���u���L���5�w|l�5~�c���x	q�O��s���&�Ćz���}l�`�I!�~���A�h�D2aƷ�b���q|��%����;"�8�,�j����~G�60+����4\�G�9h��!y�9u�5�OJ���_V�L�W<ef��+hߕZ8j>�YE�g�3a��T�MY��<�#�6�I^���Y���|���X{�5A&��W�>r��ݔ���/�;���C=���lZj��f����\���������K��HvH`Uy�H3�2.6��8��x��
&<�N!�~5'��WEWb����ZK�&C�=��#�or�UU��6�Y3�>��K֏���2�-�{/��%����i��#m$��V�)ec���i�ѻ"�ޗz��꿖��iVݤ�7z$�;�l�ҭ�h@U�W||�$�+Z+�ҜRМ�7���R�����Mz�X���팥8�x�Teni=��~<^y1g���s.w�y���c���-,���S�E���a�i1�<���S��-�����4
�1M�!��۵^�x�Ȧ0�N)}"�_\jv20vW�@�ԡ	?�Ŝs��EOI/>����L����|�ao__ns�^�����2�sCɉ5,�P����"�O�&dX'�V��M���jbu��W�3<����y�L��?I�;7���	"����Hw}�k7�����4���)ҙ21)z������|<x�d^�t i��%��͙d��"&����08J�W\9Kf�]Y����M��^}���1�R�n�U/�Q�)�c�nr�ӣJ��\����jp��t��&S�FQ���}1-/���e�lfVn�A�V�C��wVN����Un4C�X�vò�e�ƶş>�p�cbbB'"*MvE�~=��%8!��|�7�A�ª��K��C��}��bt��D�$��r ��Hf(��j��m�6�]���va���O�P�2		�b5��6o��$����c��d�φ�o�m�	Ͷ��!2~��H<��u��v@@���"6�eV�Ʋ~�ͽYd�2�b�v���p�e�Ì<�fvs�J��^��dǚs����,���ʄ�/��?�� 9����'M��T�� w)La��}��2��_e�F)�hl�PF�����,�H��A^A��p��h�߳$k'��T��`��T��A��]�3C�W�~��D��F�ʭꮼ�0/8�v���T�
?������+�[�ћ����m[�e`�z�;|�]�)5�n����s�SJ�K�χ�k�t�8��E؉f��B��#��n&�nhڈ^�4ˇ����l�r��Z��u���%N�E�&E	���`+��w�ݞ1��k&��&?i�v����B��>���*ZY`���7�Fo�3k.O���|�����?�+bK�����ё�&�:�u��]jm�ƷgcӼ��C.�f#(	�s �����)��H�N��l	8��������۞k��x�wkA�ڽ�{}�7��n�3։�Ke��f��:��@�!�/���l������X��D��h3] kw-�d7D���Zd�pk�_��mJc�ʱ/9��e��}}}Q��(��m��Դ���9�� �T1�&����5Я9�}�rV��L���i��%���I74RaL��S�TrQ�v$�G{�` ���l9o�ډ[F#�*��M
0v`uX�E ������8T,��Ce�@4NQS����Ӄ�̰��û�K����*wf6�5�Z�(���a���>�L�=����A�q��M6ߎ�ǌ������	�9���V�8��/؛X�a����ðae�G|��+�\��+i.J�����v�4��ld��z�l��&��UW�	o�a��v���0�v:w{K���:r�y8�$gټ�~j�_����;�J�we�K�p
�_�v5�?���K��:�����}��]ծ�����_R.5�������ut�Rt�ϟ?��@��[>�U)��D&wjg����x/�@>}�J~1J����aJ>{*��U�h?�`X��1
��`��+�7~�tNju����j	�[��܍���©�r$��R�b���'u
�no��J�>IZ�=_�J��2��B�s�]
?]l�����0�������7_�Bg0y��_���ީpw�
jP��uG&ۛ^�r��=pt�� Do�7k�Q�J$�T@kE�i�Z����M�Z�~M��̋)��e��ؒ�C&m�N��of��A�TE�_���|n�����Tq�>s7NY6�t�-t�Γ.������N�j�d�5�o�N�Jz����J�Y�s��o�̃h4C�`���F������r%v�y:}��X2Ia�˫K汏��ff}�$�9fCi�a?�ۤV��_T�����
�S|gv�o�35��N鋉��7G;3�?]��	��D���"�̚*.��\�׺���;0ǫ���x�+m�D����W7���������:]L��ŏ0����]�v��A��0�}8/��@9\-�x;~��g)i^�A�������R�^@��{��'�������?��(q1�5̈́<OK��_����O�h��_�����4�ikB�ۻyll���	��(��lk�8\[K+)�a�������f� 9n	R=�L�0W��#�= �������ʥo���su�����)������Z>p�U�S+�I�4���?���V�B�bͯ�$S�KD!��50P�o�ܸQ�c�	 ���,C�'�͎n���V�~B�'#rwj-�խ�6�$1|��X��R1ػ�|��2(�sAAdr��+TL0J�
��1�ҩ�n�&ڷ�O�s����[���s}|V_�7�*7��6��Y��x�za4�9��:�����z��oL��$����p���`��FY�Pj�yo�^:�.j����˻~�~�3�H�d��T�,�D��`��ce�iH�����U4Ż����:~/Ȍ��h԰4�l�hu��wl�BZ��]����!)��V�$R6{^~:?K�4�	�p�	���T*#'G$��@rD���[N$}��\|o��uRp��[Ae%%|���c�#�x^vş��kQ� e�m䶷�Kxz6�}E��_�<��o�9ڿ${�ZV_���!�74Ľ��^i��S��j����#�Aq|n�
}&�B��9k���ZsÎ7]�j�����.q�0�t���[���?_�]x�=���?O� �N��].�긝�&J��t�;;'R���������� I$C�4E��I]f����?{PA 66�r�)fp;p�;6&f7�^#�����4?���z�4rjkk�8Ɔ���5I��ٜj �� `�r���iE�y�p J��Y
�p��
U�j��;�[bl��(���X��L�g���U�� H���**1����������_��P�j[qUW�0~�K����3�
F�+灡�q���}(
����-�˹K����]�<�%D�f��0R�#�2��B�� 1:"�ٓ���ŉ)�?G���㐕�(�g���m�������;ndʊ}NDOM-/Y����0�]eG��|!�pְ�LK����m��BKK{���A�3��篦b�܂��
�]����W}���n���n���сyi0����o�!������N���Z�*121��8q4����q��Y�e���i�V@UUU�� �L'�"���r��:�PN���ae@FLL��;�]���LWm�$'J�#����ģ��d���Y7�Km���5��_٨i (��%`�B����ɤP�T�n
�X�Σߵ��1:����B�����A]���m���%�o�7
�=ޞ�������=�)������/ �#&.n;���\Y8!���BN��	x�؎"C22�ɗ(����l]�}�l�&�m =T��TJqy�q��_3�����Mٓ��o.��eJ�Q�d��{*��l)��{�XH"Lb�1�1,�c�����o�ʃ�DE�2wL�� >| i	T���.����%`��o�HO�8{Of~G^�VMK�����à۸-q����;C��?��Af�����:_�/��c?���5�ى,�G�!�lڅ�tRl1�
�CHE��$�Oң��v\i�}�.����)M7��a�H}T�:��۬�s�%y}� ��1����~	=�L436>ceWz����i
q���y��SY��� !)9"K�������S���%������%�O&aP�ҤI�ۢ=�B[@��B��Df���]���<Ѿ��gg�ϧ�!����Y;0?>��P�O(����	�3ɕl0uD��1���~�s�ۡ�ah�%ٛ2�v���{8�	Ƀ����EEत$�Ң��q�q�'m�MJ�q
����i����G~((��T���B��?[ރ�L�M>�~.��±洬l���$,����ӌ��8�βY]����d(��=?$,��8�l�K���)�?'c���QoF:f��F����`��~'��J� ݹ���ւ�̴B�A���Xt�kY�l��M.��E��*?ĹNiʊ�O��c�w�ҿ�<�t�(�%a�M��!��+{A鲴���c�t�1�(��͓O��X$zAII\pppd0��J�E�h�,e$���j;�#�L�8��j�d�
�T)��9Z�; ��zb$IO�#'M4����7f�s�)�۾'�+������d1��@D�=��J��D}��a�C�/ O�F/�ݴ�-����WSL|��s�&!!xc�D�9�����sr����?�,�14��\s׊�E�_g �� �,���V�ȟ�����<�$��YJJS�`�Q'��	���T�[��}��io�΃�P2b|ĳr�K���Q%��P1�3g'�{2d5�zj�YRJ��f�sN���Dt�yC�����m^��?�v&m ��N�֣eB���D�wL��һ�9D���#vf�f�de�:(���$s�aTˍ�H�#�Ic�wr��W|$=�y�@Q2��d|!����������}��݁�� 9����"�"�j��|pD�څbPn<�6x�f{&��D3��(7�ȸ�ԏaE���������ڤ ��n+a��q�h�Τ�<i.[b����)Ʈx�����VAq���R�J�w� ��4�/-�����нXxm�������û��1��{�'�R��jj����C�����j{[އ�RJ�������!8��Zܡ�
E
ww/P�wnł���o��{���/��X�df�<�<3�w�+��&���a)�����YO2k��p��?6���`Т��lH!)�����VnYʜQ��*tP���������%:����NS8O{$��Ƽ-H����c��������*N	�螸Ra� <�c����x���=�����{u��W��MD�g\���	Dhn�u�)ַ�ŉ	�Toog5���d�}�����eag��-k�N�?\{�t@�����4y�z ��x��l��k��1��օ�6N��|�8�7)��Ї:���G�jA_�p��= ؒsɳ��⡈����'ɂ_1�(2��ly[�\i�7+m||<6)i����u��y�C	�^�	8w��������<�B���Q{���2!��wn�0�e]*[:%*#����'k��GUK�Y:����w�e���
��A(����>���RAE38g���+�S/Ƿ��㯖�[�ra�ۅ2nd�>B�����1a��10����+�ڏ�֍?�R�kW;'���jW�A;�4jL���?�G6988�xS��Qdb��1���az$�^�)�]�;��lp��&v361�p���33��#�k՛�ϓ�ݡz�w�oq���!z.7",'��ɟ_X4��ঽ/�-�� n��V0�W��\S����;Z5x��>����:���hh3m��
�;"h���!y
$�j���@�:}ɠ�J�X���4cՐ���W�s�ϜR�io\7JM�h�L.뇶�$#�{�jog����p��裇|�8�$=ؐ����@Iz)s)u��`��ɍ��v��T����2kS[��^�&��a�V��7�CH#
�q T����Oo��X�7�xN�ȯ��+F�蟦�+�nmM�XݳQ�#�L!��R�_�'�:������gӨ��fW�W��}o�$n��ש�Ǚ3���f*[Ka����>�/�5f�r�̝)�����y�w�� ��Ps4�&�b�3��wY	�Ə8�ן'\��f_�Έ)�)��y��С �E>�����p�2�{{{_#cP2��I�D��?��Q|���tp QΉ�Q� m��;��"���p�Uc֜AM���c����A�s{�zn�;���
��q��q�a��Z��Er���f�:�c��l
�+cF��MMԝi�jQ_.TU�����`W��FJ}B��ঽ���w�����nG��U[7����|��E�WgG���$פ"K��me���yE�(X�P 칥��	8<^�����B��Urw)�-RX1P>nF��7�8���^b\�.6�S�Z���=��Lc�g��_oNx~��������r{�k��F�a	��nե��JP���<22�� �)�W�.�)���L6+bDi��nLϿ'��M� -���6�o�`_->P�Ou�5�,`�TL���8
#����_��mc��靬9�����z��sO�h�c|Ӵ�`<Խy�=st�%ѐ��]����6���2��V�|��B��7�� �%�g(���q��몿^9Y�M�e���Y)��[�1`	�f�W�p�s��w�K6��/�W/��n�6�[~�|�;�s��m3�=W]o��x�'r>�$""�3�C1�&0��'��d�:3�k�D�Z���K)��aA�* hy~����G����������������}�4O�#�;2��x=���Oݾ|�w�����7�\WSᔎ3�)�'�:y�e~h���jX@q��O9g���T*ɑ3hj�Dv�U!k$�o�ա�KOI��5 ���?�]V�h�鶯�S���-��42*����	[¿=)Kqu��1���MQ��[{��qXj�
�i�M_ўGw�aE�Z�����;K�un���(x�γ�>�`>~�V�)�q�Θ���;�� �o@�^�5I��\1wC�o�#�bM�g߭�4�Y����1<��R����W�_q��1W]�e������5��;-��t�W!2��� EK:��EHcNJ50Ή�r�j��·�p�������'�
��`+�}�w��r�u��,3�<�� ������/��'�A�6s2IG�(v���Q��a@��
�?��;�Q�R��W����U�P?�����I+� �
��"L!B	��A��sdj��k�Ù&�OE6��C����cf���D
��2؍�tJ��ƾy���q��B�q���,
��V�n�Gu�DRJ�@Ih����t-�>��J�M�y����A��mx#z�ݟHvYs�NsGO&|��!PE:ݼ`�^y�b��]M���uʌ(v��q���
���+h�+�+%���S��߆�yb&���:��_�4L�5��*�5��)��Q���^H�45�a7�'{�	��޸��5F�2i�(����|���B�t��W��
���+��sQ��xD�G�#�c"�Xӡ*=���W �����R���L�bql�0��-Pߙe��|c6�U��^D��AT{~s9pg�kJ@$F�*�ϯ���	�}CB��Q.c�~7N�-ȄX�.�h�h�Y_��� %�m�=m\?w��逰%fXﺌ�^:�pu���p���+���Zb<䏳�Ĩ����9�갊ݹ��1���b�wӄ������X/I���6ԛ�C�yL��-�dMv�����p|z�6��?��d���6��$vz
tM�K�]��F��0�eW8�F�Ȓ�ZU��/��z�N/����˱2ԍ녙F.�	��:~X�Y��+^�gM���U4]r<��qS��N@���*�����߱�^�b6:3-2u`m��Q>b8K'�k3W�>�.��}w�;k��}��Xδd��v�!�Q;��LpgW{�E�)���\Ť��8�i1rrr�I�k|v����r�ۻ����ϰ)1cUq`�!te�?Q�_��k�˥w����� �-����m������t��g���T�8��m�"�O����I0�
��k�L�FiY���R�9�;��=>�DC�N!��0U�H7�퇨Ža �:�2��E2w�'�e	~�lҏ]�El��C��,���x�&��s�Ro�WhTL�)cd�AŞ�{�@����]��D6�s��\�Hi�^���2kA[�������*�&{Hm�;�G��k���9����vQ��0i���r|2L�A�.� [AIROO�:���ahG�P0��8��#rLE9�����\u�W�P�ԫt�硝�7���<���h�q�>ۙ�5*`�*ָ��#K̐��3�ǔ���35^7o�e��Շ���ҶC8�Ka&E��	�"���h��U���?:Z���J���,{�O�����]I���T���/+�Q�bU���/���.�|��"�z�$�S��m�tQ]�T|��B�"kJӔױ��x�6g�����%1����S��\���Vu�:҃g�+�N�ǿ	� ���<w-���6��y����d-��M���4I`=2�h��>�+���!��ϟT]��x���oO^��U��8�⻷ ���ahY˞��VU�UA�N7�/�ՊM�N����+h�2���� ?@�u�¤P��uj&,�ŷ�yӟ�Mu9p���*�p�nH��+L�l7�yV��O��jc-�mێ~�9�Hֿ���%�;~q$޿;�m����b�s�;������F��n��wz��A�h�-���M�3v��pU��r�mj�N�ʁt�d�$���`}����#3~�V@�Ύ�R��u���|PO�9���`t�~���$��&8l�{�q7	���D�>�h�BxA�B��|��>4��+�<�?�����]M��d��t����)-��2$r

* ɞ@cd46]"+l�}�pr�_��%�L���o��+((8$���?��""Af���vS��o���rt�7��:J�N"��5�rr}:�T��X������v;�ՠ�3d���wNu�&�\�/��ԫ{S_�x�q�x�o�2�nΟ��uq�h�&�d=�(�i�C��(�AJC���������i#���[���Ư�H���]{Zv�Х7cw��to���q8��B��==Y|7=+�{��z��5x�+��pS�d��,�'z�2�o��C=����c��8O�Up2x�� ��A|$����ǂ�g��TX��	3.���g��H3{�zW/���~�oZ�7��qz�XlPd�� k�qv+�u��OR�Dd;��r��������u*��՘U���<9�1M�T�S�!�(�FmҧX��鶆�Y���=I��,%�Y+u�5�!YB��M.� �4�l�Z��\��g_���-졙�ˆ�֥M�N&�������b����䣌��L��"���?�ɱ��V�\Y�ԇ�P�<���I2����nS+�V����k�����ml׍�A@��x��E�a��F�j����~�ǌ�����.ǂʣ[� �A��j���.b(�.�3.�5��pޤ�\��'�i�oj<��,~P�Nߦ�ǫ���b��⳥6�^�ZK����F�a�p{�� ��g̈���԰a��C�2:N�"���_��YA4$�63~���g$��d���r����̦�Zt���j�%�ν��V�������t�B����@gX1p",����Q�s���1?m@����~��)Y��'��t0��I0�n漭Ĕp7u9�K���W�\Ϫ��vC�i����Τ����5P�n�U�'l �+�ö�����VOO��A�\U ��B.~a$7m���E2b�q�7��,Ch�ފ�I�i���<�"^�	NH�(���]zG�Ǎ\۟R6��H�W���6Y""<�g��k�A|0"�â��%��������6t
|
��X8L�K��x��`�K�\��ϻF}�M^��Ґ>6����=f�و"K�͸�(�ok�\A��Y�nu2ݮ�D��Y���4�=�9;Si���|B��܇S��<ʀ��n���;iᓭ���Q�]h*���,�$��;�*iʺ	�a�t�F:W�h�S�ڸ�Sp27����8��
�!kY��|2D?�,����t�������c�In�b���aX�'Ϻ��c��8L>�[����L��F��� <k��f��r��˶�T��8uT����d�dB�	" �C�>a2TW#���a��Y�#q�a3�V��r(��2��n�  rZ�:���  v!��Y<
�\��yA��@ʡn��"��1���i����0ӈ���.�,����(�Y���y�B����F'e��T������Vq��utQ�~J�]�#��yY�@	�����9I��m]�H�*��ŉ���j ?��i��Q���H/��M�!lvng�)93i��gdóJ�hy�vű�L�T�!@�1��$>��X(Ք�6���y%�Ô��w�yw~�w<r���b�=��H9���X-���M��.��.@A� �����z"�� yyޣ]��*�t���J2�8�Y3Ǘ-$�|"����>DN�@�Z˯`�ڭ`����E_Zg>|�u�-����=ͷ��:2g�=t���,�/SnA�K��b�%.�>VI���~=����Z��rh�4�0���j`6�s�u?&�?��ؽ�Ƽ�R>l?މk�Iq���z��4��P\ا�z��=E�G�Y���u����i��qsr�+���}�J���F�N�\W��f�7`� {��PJ���op^`E�+D<4�_����k�"��=d���������+>%<�E�)� 6#c�㰟D!N"��G"p]��ř;��Ε;ٌ7�*�z���1���?�-��V0��ַ�c��8D:{r-nV�q͘�E����OFĒ���ら�E��#ĩ1<������Z.,N����vvwc��^��q�'{U(u�5�A ���	-�5E2"̖(c�#e��D�-���2m�����r�N�	� �uB�0�'������DfT}��z=}�ð��(�����=s�똏ݐ��AV,�_e�?�l��p��V�,g�to��io74�>���_k�_��~���x���:o��t��5���t5wg����z�a3A��XlI�R�͈''/�R8�,	�V�3�Z��+�U'E��ϿB�#즎�R���Φ�+��-�Lה�h׍���#��z�O�.o��z�L���~iH�g3v?AWl��nIlΎA� J��%�+�ԚS�b9��vBH�!Ii�<V,K���5��z)r�~z�W�g�����7VC���R����~W��ǕB�.�Ϣ�p���1�qt�D�T�Ӏ�_#>=���j��ԙ��Y������MWVI	�U��#��d#�r��JV�IRҞ�c!^Js���`z��w�ݓ�_�rg��b9!/xѠ��C�-�.��r�Õ��Js�?O��Z�����T�:'8� ?�^�n��uc��K	ё*�Ҿ�6�ÛP�@��k@��v����
� l�͛��v� �]�_l9H���!���7���#�,�[5��()�T������UD�p ����q4n�I�@���:Z����?>0�2��2^Df�	zK�y�� �v��.Ru:e���R��߽����M>u�ǵe	��g�H�4cMs���${���%J�6jݵ�ݤ��7��������'����2^���o��Ig;�dYp�X���I�әN ���H<U���^��pL��A�K�z'%٘�3lYD��E^����H~�b�����u��7�fe��ڕ���D�qF�����I���l������9��)ԉ����h{�2O��&ӆTh����N�4���+�()tTG=�S�,�5�wq����;,��˯��Exw���n�mx������sӬ�4x)�]�OT;!���%�)`�r}
H�f����lc-���U��ܼ��Ԇ�<0����ϓ:�5/#���t�6o�
�nF�;RSr'WL����]e�֤<��B^�h'gD}�'"��L��N�ԛn�W&���~�\���|CF}�X����?�N�C��׆��d��U��A�R~/ñ5B��u�xzz��£dß������b�f�>d=5�]�Ƶr9q��_{H�Ӓ��{��D�j����w�|M`�r���L�s虨��n]G�bj��w�PAF��ǊJ���#vu�_�c�#�]g����vM|��I�+0�T��ރ���sB%u%����x�iԿ��DP�&e�w��\y��ɷ,ג��x%(�&&��.�t��2(S�<����o
�}� �� kk9 �7E֖ϗ��q�*Sc��!�L�a���9�2�.�ʏ}�;۹��S��3���g�F[y��}�A�G������`�0�lSݘ�RI��}ѩ��"��uM�jjb��U;�jQz.ꩨ�E��'�Ŕ���	/�V�C�Ez����N�#mF�);}����k��<�'�7}}��Z�8�UTTl����O���q�'*��>��?���%ì��-.��Z ����r��z��{�3AE}/���h��_
�y��&5���on��AhZJ�@$b�x ��^�Ձ���b	X6M��b�����o�]P$~2���B��C�a����Hl5~�a7�e�B>��xO�KcZd.�wDZ�k���v��$�(Z`l(�_��o-��<m-RBXC�Z?�T�w�C��G=���D�rd�R;��(=:��IbY&�M���V���H�W�=#=�����j!d| [��j>���m�N�,��}}w�c �Ӡ,p��\<�����������'����e
����@eJ��}�xFԻ{�	���ä$rƋ>Jd�̈M��������!"*J��Ptk���4v����{DN��W��Rh1Y�Yn?�5�qi��fq�ޖ�7�zz6�6	D2| �ui����L��N WU��"0����(��Ev���h����,���4c�0/?�u?�ˇ������Yʐ�ҙP0��V[��z�m���߄��K@.k���G9;�ۮ�>�m�$agR�.&�-� g}i�33�Z�N&��e���@���޽ �[�w�E�����ׇ���Oc�G,%�h�0��\7?�?�K�M*Ot�l�?��ʑ�����k��=�lpr��W�}||"�X�������W>�[����.t�����+WE	A�׉��=<x���p
vo�e����y�����l��������� +͋� ��'�f0�_(^��Ur�O!�'���%�lQ��#�~nj{k�/:��!�Sȸ�=�q�E��:g"wN|&�w�q�g(eK����C��{Tb�y��$'Τ���}�1wN�\4����(�u"�l��pC�mHB�@Ț�E�k����2��,�1@�M����`�� ��	�cy�0�c��yd�F�Ic�Z3�ؠ�kL�[0�w����E`��Q�m���W.!�����J���|n���*�$�cC΢Sm�:��Vq�U�y[�䌿"�z���b/�
x�e�T1U�!p���Ȓ��'�ΒI��������*��E�q��1��iٹ��f�y+AKK�H'!���:����r���]�B�R��ץ����}.��W��l��
�l�a��i�ɨbyQ67���i�\��q��E�"��䭭���#������NӸӧ�}�X��g<d=3\���s��B^�Aß�g b7����|��O_*O�ٰ((%f���5�V�ѦQ�sZ�]J�{~�!�XO)E�vX-"��q(��0�֬�+N�����[��v�1����6NoW���hT��N�`��!�+���nʢT�}mn,��.7��J���yޣ}�K�!t�	���a�����+2ti��?��ъO��ƌ�'�cG�Y}�ǟ��
�&᰷�S<V����
y'�6��g�{���j#�������G��xG'�Qw�5��i�w_��ӵ?�'� _Ў�畔���&6g͵��5Wyd����"l�:��:3��G!����������H!��,�~8����Z�4�)3�u��Vފ��� U�v����vQDd�� ���{*��E�%�Ћ3|�q�B\�AR�a)m!�z���R�0ų8�xm�0���F^�����z$'k�-����ץ4z�NwM{M�D���H^_�X�8�r]�	BCc�[���^�+�G�q��?b���,E �[�2������iTϵl��ͬa�ƭ.ט�[�x(~�9�
�w�N����c7�	����b��>JY_��&�|H6rv�1��#�KW�{�>�_�M*`�A����'�J���{b۶jĭ��2Vʂ���k��^y":���H�.�a����۾�or��A�'�W&��U�.q�{�� <i�G�G� pA�����7f+�LNm��BQ���J���P�"���T��K\;�V]���"Z%��4U�-j��?M��*E��5;�>4��h.0;0n���M�P|��.v��L�M)�o�w��������L��������J�^XaKTj�"�n<����[�X봸`�(�EKeOP9���\s�8~��<�����������4�o��?q�uNwe{�� q��g[�Z�=��>sΨ:�u���\�x���o���|�G� ƾ��┕m�)�Ζָ�c��.uA���vB)*�%z6p��޾����b)+b#I�lfBLo�~oc�{�D�8�P��<��Ğdn�e������r�!�~�em�7�!����ό�22���I/Ձ��`�]I֎4��:���1ɢ"N\��gj$�
��E|��H�;r�n
�]9�_�j��O�)N�OB��Q�ϻU%�����U���g�x��%b�x�d$R����1���'4ZtY�����ן��ܱ~45�	V/�)RƌM�[Z[�ٹ�O%j#�y�^ڶ��w���AO����n�\�ֻe8��Z��
�'T�iz���&H�W��QF���;��F��QT�\��]���oW�s��LĿ����v��̝U���$�7�B�+�D�O��L�Z|����wO���Ş�ٜ/�]UG�p,'�2>�^�M�omT4��lY)#���e��_��3(���f�G��;H��V���f ̪N􅁊��
o������x'�V!��?Id�����~T%Q6<���L��^�%�=V*���a߆��7;;�?�m|jp�:�^&�ζ�ެ��"��l�	�"aXe��i�h�=�o�l�N��E����m撷��$&��:g�}�a�.K���ZZ�z�^�;��ҕ�	�Żkw&����iłt�O$�\[]�t3���a s�Ǵ0���Θ0WB�[�d����U���&�n<�+ז�p�[�0�+���DR�l�I��t=|#L#� O���E/�
��-'?MBj0\��Ǵɣ�E����D�����Q�?�����}�Td�^pBdHua�R��ˢ;��_�����g*/�yT��*Z�[]�2[��aֈ�q'����(����bnR\��R���:0;<��jx��v_CW=m?V=�����"?A�%Ǻ��d�4궠^{nn�����Q���_�	������XD���"��t!�%��L�
&��<�'"(H��S zK{{%YY��GX��$pi��F��:ٛ,�t�Ϟ���ƴoq�Q�s�����)R�))����P�HK���x��i���CT�(l��*��v�e�@`-xq� (����ͪ��L�+�G�q#n����� �[F١K	UYto�W;��n
����%7�k���O2*���#�d:MBb���:��؍��~������r�;�n<��aG����U�J�׳Ԙ�:\Y�x���w�=�����[�?�^�.ʞ߈t��o�:�<2��'�}�GzK�F�X��`%r0�|T���  ϵV�R�#Ǝ���z�j�1Z�����)*�3s�t��&���o&v�G�������KO�hu|���7�P��T]�Sj��0>�M!$��������a�1�?Ѿ�RZ7� ��^eF!�y)Ƿ������5�L��u&�~�������ǃ�	̨���b�з7�H�u%eD˷���-Yt�ŀ�P�����$]�7g$��FT�ڊ�̖��c��l���N����~.��/�0�"�*�_�D�nG���AR���\ZZ��E��h���>�⦢�M�FO����2�a���ص��M�N0���_���q���+�fgm�+�[(TIho��WJ�/�L �?�<u���rG5p�	�d�U�\'��$� �l
u;�J�q�a���.���8��;�m��_Ge%T
�J/����%����0DA��B��0 �,j ��+�A�a@�#eF�ܒ��;�̩=� �FBD�����ex=*pu����$�Dp��lt^v�+??�BÝ�{1�[�R�#��EϼGDt�S��l�Y�d�0��k��VJ���Zx!��ϫ��4��Q�"P
��Msd�a����1�,�Ҿ������hQ�׵����;�d�l��N�5ip��Qsi?�?�����T$��I%������9��f���b�3y�:nC�9�;�r�
u�<��X��0i%/��k>\�뺍$F�|z��,U?�HO��-C8�nO��W��毇��g�} ��g��� ��ɥ���@�G��P$�@�T��+��S�v������h%)l�z4H�w5���N.jl9�_Tϔ[q�	\!^!��ߐD��`9J��J��-k�<q���ՕX]�S�&x���F����ީ�³�p��e�_}�#)����ʿ�D��9������n��B��8z�o� ī�$U���e+B�?�A�ɒ&���&}�Re�p�>c�3��>y��������0���7�̦�[9�^�����6��V���/��E�)ko��TF	K~i��E��J��`P�U���&쎈��k4Lx7{ޠH;��p�QA"������=��t�ǌ��sbf��f;���ǃE��v�B�4������5ho��=~��.�ij1v !�����Cl�n�����j�o �A���v���Pj]�&���Fg���(�k��&f�>�2%����� e=r	Q#�S�X��CJR��)��¿9ϳ
0?mܓJ�|W*΢&�Դ�vnix��)�r0���(b"�u�o�?����J=K[k�c�j�ޒ���9X�~k�%YU��FP#W���ݰ�������R�Y����"!!�����,><�#�E�@`nM�	�������ki�m����X�Â���+9�5��ji̢2�I���f~}���Z��M9]P�7��_�?Aj�M`��z&����c=����-���<��.%�4)��O��o��2̞*x�p������mS(����tw�o3:q�� R�'_G=�P%��Oy�pC�vio<ՍW�G�L{���G�Ö��"�M��T��c<��X�����E52�Q7�u&-w��[�����ve3W޳��3����G���yd8�^.�s��a<`��E����M*�3�1fE=�M�F��n  ��e1Sa䁶2���0J�M^�6�v�+V!_IN��U�|��n��8N1����F�}W�~�����_�z���c��>3�4����}�\��L4n�+��5t!U�#ٛ�Թ�}X�A-*`�+P�7A��}��Y�.�)�\~)��Q�̾i�˱R�!��f�-�&�U4n�,������fJJP�bW�����k��L�D��H�Y��k�3�;k%	RUsu��^��-+b���3�G�GS|�/���,`��%Š�v�:J��vO`E��J�����e �^ݦ;�pݛ!XKg=���Z�������ԕ�)2�HV���B�LG������"�����yjbG��� i�^�ڞ�:�.� lsǃ�k�\����v����iϽlW�*<s�{f�F�F-F%���T��}t[j2h��;! ϗ������G�������4����,ۧ^�,8��|�¤a#�50��;����E���VG4�_
�]��R�����ϰ�}tf�DjJ���Q7�u��p4�3S�,�p��@ ��#� ��a����m����YTX؃]�`'�VUd�q6Yc��q�7�q�a���?Q�k:�g�D�@+$�g��^pz8<��_I�P���@c�&f��I⃈ed5�ݍ�ls	;_��G󅪛�`:�� �9�E���Vހ�Y�f�歾�+�e�zTnO��f�Bu�8�8}��~}���-U�3m�vz��>�m"_~�]!݄��a�g-@` 1�B@�E���K��YbÈo�&/*��ޑ�ϭ�oKh��$zQmc�5�!���%��I4x��E���'&�q{@���;��^i<���tЬ��X2�z�7�,+�&�������H�M�A�$1}#AUK1�W�+
T�:'�s�� b�ي���#n%�5���(.�-[
����b�����)��{=�R>��
����VXIh�(޺���Y��h���-N<w��H����m�a7����?9#���R"�&]_�:��)#�e[�kb﨤���)ss��x�%g2c���V΅���_I�gΡ��QcI	�����=uA]�^����-��y�U8���Q۟��V�'O�6�>緰$0X��8��S$�~_�{@��<�C��"� �n&�p�.����m!���899���s�nV����'_���h0�ޠ�YC��C?���"+�lH�&��U��`pڝ���B[v�B[���Wլ#]D4/3̥^�/��22=y�� ��@+��~U��8wc�P��~-q\{�k{�X}J�<|�繄]�K82��ej��Sp�Q'�7Fh�����gnY�)XƷ�Mı���j����M�sW"�&����V�6.��iX[���*/�{�-��_E�5�){������6
V��D��_����M���5�_�HP���a-��_A�����������:xy�8
�1pe�G0D�����p�e����j�g%]�Ϭ.��#������̯GF�ާ#��m���,2�)RG�2Pd[%�O�x�� ��F�g������'���dc����d|��+t�P����ё���`aNN�݂�
�҄��xך�*��(�yAJ�˄3��	3?�$�H�_A_O���v��d��\1a�5��'�m���f%����T�C2e@n��d$��S���aWg9�K���G�d~TqY"z�4<Jz8}��\i�#����Ë#3��L ���J{?J����fV��\�Q����e���+7d�몦bKA�͢��)�G�{�8���exܽ�c�����ߧ���T߀0WYb5a1�.R�{��Y���e*/={��>�n��W����:9\+�UX֛�����6b���)O�9�$M�(KcI�_���Nz��ޡ�a(��%���r��E��@حIK�?v�-�k��e[����}��Ǒ��3+���ު>t��sjW�3��D���S�'��H� f�|����4"A�W�̸q���,�E��B�	��hss�����S�Ö�/�Q�y�v߭Lk���z]w���Hy�[�v�r�<����=m[�b^�b����4�ߧ��� ���6\��M�q�X���fz�l�x�p�ۑ���P0��P4d�E�n�`kf��
����G���������K2���3�L��O�;L����R�q%�|%\{e{f~��O�:�cg��h�`��	C�"���B�do�#9��?�����J:�r���2f����~�ʧ�;|�݆�k]-�A��O�Vĝ���t���w�m��)�$�E|ϕ,��J��5�_��)�L����gP���v���l�.�z!/���h�k��w�	�P$�o6M��"W_WYXvK�t0_稐ix��ȔAUyT$�=�V^l0�ֵ��u� ��wΠzn�EpP�w�!�*�K����s�=5���a�n�I�:G��%�/c�,�ܾnI���(`���{h������f{&{"������1�0�/����D��	�=���]@��� 4�&H7ߟ�^x�N�-��+hnz'g�R��n�P+}���	�o�ѧ���O��u�����a�bo��5RQ7+KQ�_���x+M�La"�i�������?���vD����e�bh���d
?���@���ڭք�ߛ��0�8��,P��W\��wTH5�g~�/�)Zz����3C�o�-��1a`�ҧ��x?��O�	;ZO�=JG��<wP��9��4��gP��J��R/�1����{��e�+�^�N�{�'��O�e����0�-���{�(+չ	?}x������Y*��+��z�e�9P�t�RN5Q��k(��⬟�������v.F�h��ň`�a���� ��U� xT^�����*�����`
aR�,�n�h^8�H7����/}����(����4ī�%���W�d��1w�-Ƞ.ɵ5�z�7�}.1[\�gM���W��ˤ�����;y�Cֲn4V�~_5[�+�HIo� �b�K&����kr��-C��xա��U&m2�FF�bE�J_��c��2�|!֣E�*O�8����u��a�3\.����((,T�-[J������(���8I]�q���DUJ��������d���扆J������f���u5�)����}U�Z��V��чt���L�d��6�s�"�V���'�<���v��YDp�oEѿrP�o��ˈ����K\�.�ʒ\e�HO���e:�JF�>�l�tX���Eg\���K��)���r���hK�`�W�^-���� ��������z|�(lRZ�)��,}�	Y����gĹ�+#���!~s���ᓠ���6��K5޳��ffo�j=z�E���p"�b键�s�ŕ����$����g2!�e��_���1!�>��>_�%�+.,,<�wП�B�������>>�1��+{6�hۧÌ�p�?u�|Ѝ�Ho�ꍸ�H\w@�ȧ�	�6>K��|^�j�������[!o��Dqh᲎����t���v2�~F�{xs�v��k��%p�:PW��
!m/.`_oXS�a�~	� ^�Xߚ��gϋ7���Ԅ������x��۾y��Zk�S4�0c��8P=���Z2��]S��H s45�X�V����H\+̥&�'����!^A�R��0�r��cU
ITE2�����&u*�-v�F�y*��*2`?�L�Y� 7��V|CS!<IUk5��68�F%4L��lG�۷���'	����6��O���:��<x�u���g܏]6���=/���,��"�:C��	߱��Lڋ�lNu�"�?�d���`7�L�M��j���,���@�{�<��3��'|edaR��[0g�W��c z�a�H��VI�8yu4?���j���q��#���ց�
��su1���o�&)�v�������>Sc���O=��>�f��٣E*�uI@���G
D���,Am5�4B���L*�?���d��h����}���VZ��[�%G�c]�i�U/ѯ}���6�/ >�e�0���9Ҡ${�W�1#x���TǪV�@�5��GU������e���}ϖ�ዓ�9$]:7�-d�#��;uc�=>��u��]C�jV�[N�<�ԝ �P�H����϶SKK,0�7by�k�yhO�[�,�gh��BQ�ѽ��Qt9�u8F��7Z����)�SPsO����mk+�S<�;��E�������iQǘߌ�o(R�o�g,ԍp ��M���H k�������kK"�ZnC�4�Dw��Q�l�B���K��F�R�3�\������,*`�׵Y��+1\�4����D�3�΀��2M�Y!^����ͣ�=֠��l���Fz�l�ݳ\V��ս�����`.�i���<��1�T=�'��dk��bظ���r'�X��3�gfDT�m���-S_�x����ǜ�t� ~�6����2�m�P�ʕ��}����������  ��瀇�	�����[�E�=�ò.JH#-��]
��% �K�(�tIwww+��H
(�y/~?�����G<���3q]3sf�,`���U��L!V�S�U�^lv�SE�&Zf��ط�nc�`�� s��H�WLYbӒ;�}̊5�s��S�4 ���Cf
��Y�T����ϭj�A]��-J��P�cQ��C^�li|�
��Ra1����#r�^������֭*�ww.e���ʛ�TԾ.2m)"L_�6ӤhM�Ԝr�.Q�����7KRhn��4�j{�{	'U;`mX�p:�����5eZB�73����(E��F	����BBB���,�7�;[[!��<��ld��8O|_r��R;+&��F����(n�l;�tJ接x��~x��(c`��ʽ9�ׄ��&
6F�e��Й�9�dӶ���೧Um7Թ�����cu$��H�e-�懢����gժh����Z�Ko���S�l��$����E��(��F��$�ly)����/�9�ڒ��@�~>V�j!HR�;������.�CA8O)4��l�L�0��wne��2999�����d-�@1?:ӥ����]���o�w���5����%�fk����3Α���ƹ�<��G��!.�gO�%�_� �=
�ɝ�v��v��p�4�3`6^�9���M�m#�3`ʴf��n�#�IK�4>�r7Xj��N�'��J�睹��	XX)t����XM�04�ܪT@���3_r����5p6ו)�X��� �ĺ����E�v�C|Q[@]'��)��&r���1kl��d��s6U��8�U�A�BL��H��[n�qͅ
�ůe�x��s���V����7�%H���u6_ϥo��޼�0v�d�mD��]r�Q��'9S�l�*a�^����Y��'8��������P�&{�>� BrX+j[��2�HA]|_;7�bѣ�0c�df,��9/}3%�zXP �TT�$�����Sk9�4��t�v{'�F���U�����3$�%��\����kh9zˊ1C����67#��g)bȽ� �U=%�X�e��\�����������˪>��N\G_XOWf�X�z	fK�Nd�����KZ�o��>$���iͻ�� }ڡ�?�\6���Q+�˙N��Kۈ� Ʒ��߁��������9��p�bE�ǻ9=+V�nF�W��BC�VH&̪;�f��g���=y�ư^�����N��1f;�k���:I&�i2ӹ�_��h�d8��e"E���	d�X�^�J���G@.�F�b1,_I�io���̝��S��ڑ��%,����_���Unx,� �d�U�����1Dɶ���~�Z�k����'4�e���Cqb"8ưѵO��c�5�T	�ڝB��Z��s>�`�G%�6
̬��f[�-�S��,S�D��&���0�������H��Z����葃:5�����	��޻Q'�u2�{�ۣ-��R$@k 3�!�,�Q&h��
��A�%�	��:��@f����l�04�r�߅�ޘ��܍����þ�&��n���#���%s��徺��d<��m��˾�[}��ꃆ}��w�lJ��
��w��*~��߃f
�H�ҳ�Rbm�Z'�ꄟ��bVs��d��fE�k#3��{r3
�]*U�t���,�	���i�^��88����#��^�ܭ�#Y����,R��]c��"�=���eL�K< ��-���G��?n���4(�����0JaLN�̄�G�GL��^��I?����c�����M�9�N��Y:h�:h8���>�{����!cgx�'X���_ZMݚT�'�ܐxk�`K�l�!3΂��-�36l����]��Cǌ���a�T�nj���^��Վ��w|5�����	6��P�ո����i���W~^5�yw8w䰳�Ij��М�4�G�L�PGfg�?68`dr�MXP��t���'�|�R�%��=�=�d䕌dKpL�%����?�3DD3�����;e�M Q��q�	[�IkY����>�#��ƭC?�b'Kg�y�p]������l��᾽����U��t�D��c�aO��2�į������tɵ�ϔ�b;ux9�?h�Lm�L��+UZrV���������U���E�g�)��'_�0�]��P��Z�����9[����\�PdR�������B�t����,�a�Q�FQNP�궇��>��HᾸ(�4���@��sY��O�mK����J���`t|g!1��{&�p(Êq�o��`�t���_������m��� 1DM$�\�P�~�#�{2�X�T�ac���=]{�&c��8)��h�+����"�z�����^%�Z<�c�"i�����b���o�-X�����=/������qc�Rzq����܁������F�Q�3�
�r����=���̠uNV�>�4�)q�����?�Y1�`��u`������8ӸZ�~���/J�׺�ߢ���ĝ�����Y'�)E��z-Z��k��
��t�a�N�k��bN��	����Mh�����7~��w-~�-P9r@^�2�9���A�=^�N�{j�5L���E�R1H8Z?�����xm���zl�����A�+�g3�m,�E	�^�=�b�fae������*�8a�(ʳ�d?��:t���l1��C�� IE�{�y"L<N��8z�2�N�/�l��göO�N��B|�(��>�0]�%]l|z߹;#�wІ�ڕ��o�-�li�\GD@�V����0�@��l��u��N���6q������ڹŀy�Rܱ˗F�B�B���(��h̍	J������Oڋ����y�sR�;��O��9ƫ(2���OT1W����_��B~�`f�/�9ԃ�����Km#n��R�9f@���=	&������EL�Av�<9��D&� �|i���.�{5D�����Ta�o�LY���oįA�r���aB27}��`[O��nm�~��<N��j&���DTNeg��Ք���qт M�UW��L��*��ã��R!�A�$�����f3��=��A,Y�̳gO|?ﵶn$�=x.D��%��R���ᣧX�ܱ[�M�[�v\�zh�P�	���E ��{�fK�'-5ō���#�\���
��_{m�~���ں<p�+��ì<Ǉ����^��r%�n�d�|�p��j�|�U��\�$�[b�����t9�\�
���Ĉ`�G׺��z;}.´p
�{
m���CꩠZ~� ��C��Cf�9��CBB@0��YYs,��G�� 6$��)T�{*��%iI�ʭd���K�LG��
�U���t0�Y�Ɍ�t4]�;�q�*�׀p]ꩻW����1�.�_�S��&��0~�� ���O4`ŮpK��*X�������ʲg`�Q����1��Ϥr�$��|�Z�=���=�M��A�@+e�ED��1��q�� �)_�X{d�E%##H�q?%��ĹA>��F�V��MF�ԡ���l;�-��T2��QO�2���X���Ϭc�U���Ώ�&��2ܻ<�]C,�02fD���o��bs�w��^7v�=��D	NJ�*vt���]N�}���m����	 �ɸ�G�4�]��p۴�3u�&(����V8��k�$N�%����^�X��]}���JW���.�s�#`}%U����p�mS(�w�����
�����S'V�ՎZZ�4s��}�/d�>�I�2?�!�&���E����z�m#���#�!XI��ؔ���qO�}��I5Bۯy$��7���){�~D���i6�k.�K]TO3�4����j!��T��E� �2�=ĶeM�;9S�Js�?�L<RFNN���羦�{1R�������~h7..nX�Jޛ{/���  �"�����&`)4���ܺl��"!���t҄�Wu�]�;�������҅���'D��> ��ѵQIK�J����~�ۊ�3�P��甪���gπ��T��m��y0V�D�"�i�!�eˤ�!�u����Ф<JH���tF�Q����QS�ϟ�-~BP�R���d2���Ng�eW��l�6	(sZ
mkJ&\U�l�Pϵ��9c��f���u���
��3�3@��Z&��k�y�)��|=@�͚�����Ǘ�kym��N'�LPYP0~I�7@fc��I�һ�N΄6�|)�α���_:�B.�?�����(�9���t��X/Ʒ^�� qBġ}>���q��p~ڽ�P�o׬A�!�Цw_$��lM.*Nʛ�'�N4�n�ty�i�%��IHHB;)�` k>�����I�,$���6>�'	T��l��|�����Z ���׷"�6��u��.��PN �65;;�� �l�=��D�&,�{vg���D1Q��9�X9�'hB�gwZ�
��Wc��vH<�V�9��*��y�f	A�s�.�#����*�S�jIEK�cY�v(�YQN���?�9^1�sx.��������>37w�)�mU���F���S�GK�6	`��N3���նi����!�O�餉e�ݠ�x�H��k>f���X��b#Tj�� ����J��0�;%W]1K��)]���}a���O��{�sSe�����րR=N��q�L�}{�D�Ç |���3�ݿ��܇���F�����*Ձ)�� Z����^KF����n`+Zw@;#����R)�(���+�	�^��6�j�!�0�w�r��@��H��k��Q��sJs[��ϲ��Ƽպ�B��@� c�6�Л�x�g��ܟ��)���&��p�{
���E�t>Q��&^I�57���3pHf�J@l�/ѿ����}�*� �P���ABƃ@|�v094���+V�&A���+�q)��"#o��R��L^�n����i�;�v�|0,�,"Hq���(��v�\�<)���7���L#g}�ȝ�#]�����1	<-���w�8(�9Ce����jao�xm��8�lzm��ǒ��B��eB|��N���Lf�V&7�`���a{7�`��$錫oi�{�i��}i,���1�W�p�t�粁_}��^@��ˏ|+h��t����<���_��V0r���(A��>��$�B�cybe�e�����I�ZG��)�"�Y)��K]۩9Q��O�՜�~�!���q��Յ�� �zV G�U1STxH��,���u�<�aS	54gSvR�G�"4+�Q[���X�P璬Gy�����Ҩ���efx�+ӑ&@%�F����2�)���n2�1m��^�"�ބ���`�z�Tm�*��U@�X�d�Q�^Q���Ԯ��{C
�?�z��^BfW%(��k�w'�;�:�O�U�$�߸y�Y�!�w1�`5T�-���t�A���2�&p%"��ٗ�t�&�C�4�oj60U
�[*#�]7`jQOOkH���O��j#�δY���46O��-��hkF�5���6H��p�۳7��R1��'��O炨Q��R�91J#M�IF`z���~�K,�7�%��x��)��\�`�Qr�_W��(���kԘ�#�͛75�^�tia�C�c�7a��KFI��� j���C�@('�����(p��%��o�g֭��&�mP�]{O��P7�y{qpp�i��O�?�'�g��1ܜ,qI�5�섛�,���X���!�Jd�9�@���O~7r����i�U���l{�ø����Z��襛]�d��|����t�_�W�<u�!�I)5;�]!ݝ��%u;!v�4²��^�(������|��`��W#�Ll)�8��^_Q#&�_O�x����]1j�#\�J��<ߍ�,|��~��r�=�7��e6���r�K�WY�W��Ѫ84��!�a���O֯���#�3���U���Q7Mm��	 �����1���j >�o��K������ʭ���.=����݈�%�Vt P���^��r��V�_X��vJ[�-g�z'�^Y�W�6��5��<ק׽�>"6-��,e�@�b�C���t��C�,B�XAG@�*��I�0�i1=�)�f���s�ý6���q�������IV;�z;H��f��j��s�~K� UZx�κ�1*iw�*�D�K��.F�t|0�����C&�����/z*mTҮ��4�ܖN�#ח��C4�2�֥���L���E�Q!H��a�)Sh �ˡVz�T�=�<2�	�����J�~7"���T��k����<���s:��^�!6J�n�(��As��⮕z���*<�z�.h ��L��_�-O0�͈ª�XE�Ӓ�jDٕ�P*J�����h�|Wh��h@�g�<���;+N����4���4����G�Q4iB�7�ɛ1V�a���h�p�t\����h�H:Z�p5fu���%���~��D\�J��QɆ\��7�%<>X�_<���l'G�w�Qq	O������_�� tAly�]W����O����~�Ģ��|����qp)y`ً�u]���3'�.����eq}Oxo'ۂ�������H	���S�Q/�l	u�v�NT)m��)���҃6��x�����biG�z]�8F�{�������Y���`[��HV����ێ���67��Yw�n�$�鴾��C�i�r�}�7Djn>'�&��Vy
�}��>��'����5���+,�(H�#�F�/��R0u�����q�"��΄�R%���v.�W1\��E�-�f�A�,<4 *ȚTgF}��<@R��P�̖u�0\N�f,��wި��ֳ��3���c[U����fVV*b�Ջn�+͢�QF2��nI����jw�� �$����}4�*y�K���7E���f�"�A���Qn0�$�Z�k�1�#���^NG��rU�F�_5x��V ���4���?<���}�3�/He9<��T���ỳl�b�u�3D�|��7/Y0����^��)������[�'�Yk�C�uuGk�\��ܶB,�߉0��``s�Ka��)�b���Ƀ��PP��Q|����zb�u���v�U�P�T���[���h 5X�p���4t�c7qy���
�T�:}��?���LOR������fkN�����k��Z��E6��!�\�Y(�Sb�f~M�<�'�o��t},������ǻCz���ǔ�t{�c�+�/j�m�*�À�-D��+�>Z��c%�{�j}��r!����l�ި�8��D���;�:aA�y�?���7��A2y�/%�;0b`�X&9E�=f
0��`wHY�Y�S���������'��MOQ�}c���h$�佉+)��ۨ������L���:�yc�d�˜$\*j�S���q����HW��{�����{���So��Kt�.ƅ���"a"�%.;NH���ny��E�l�c�O��R�=*W��
��1�>*�;a�E�@��w)��7����4�ѿC,���f�j!R�.��ݓ̹�[c���v�Hɩm$ex�ʛ_�¦	�{(=v��27��r�I��.�VQ؇g^��� a����~��uT:��ѹRj\^���
Q��6�����nQ��C�n�Ol[����ƚ~�VT��ҿ���
��ŝ;�-�3�kvu��;2���e,hm�fK�"(�-��^��ӄq�9�ǿx�% B���+E���N���1�}~����.��Tg�yL@i�la�m������������z��g��7/�Q�K���V�m�h$:>ܑg�8�6�<h�U����\�������Gޤ�F=����t&�$E�S�3�义ɲ���>�!��DK8��!�����l�{��qc�3
 �����x��nA4���Ǭ�f@%�����u��V���`��Z��XZ*?~l$W��6;7G!	��-U|��A�P������xL}8ABg��-nW$ NQA����A���/ֻ����� 6i�J���j ��F�?�jң���xm��j3������L
��noи�Ͽ��Ѥ� �q�/KQ�Q���6���8G���^C�>B�]��>Ńd`�IIIQ���=[�u�@��($#�=�`��I�L.]�75�X��G�����R1�	��2��K��y[5Z������6�h��W��f�E���~��d�~����ݽb�7��34�cB<¹��Ij+�3�V��͘T�K���e�'�}_��o{�6؝�yx�������Xb������󼹫�<���������&&��,^��ڇ�m�1����]�K�\C�����6��r韧�KR�V=�j�a����FBd�����!��׎���ZY��(D<HHH0�>!��qf�wp�k��F��e,9_�-a�E,���o�2=��*9�p+ɼ�����	Vp|R�ꯈw& �ߍW#��ot�1O;�n��K�����е�}����}lg�I��������!ψ��(=�2�]��Ơ���ni[n,�zU���q�ґ�t�l�c��"!?���-�j�P�gJ�9�A��)	m���������.�YMƚ.w�K��f��dۂ)�}Z�ٷ���;t'*�I�H�+��Dcm������俦�_O`3��H�,��!~u��c�k�2� �K�[�8Zt}/�Ec���ݡ?錓Chϰ�k��^��_�o%�����z���cWI����x����|}j�W_Q��HL
F��&z��Ɔl�E�&�-#&������ ��} ��{�] ��k��,m08ߒB� T�Y9�|�c�vd�uL�[��_eb��|�x%��:��z#_�i~~������X��m�rI������[��_~	Ƃ����\��)�k����ro�]U�)ŗkWQ��\u�������^�<�K�ϵ�����}�E�>}�� ~v$r���mdo0Y_�&�N�_�0���4�ŘH���SpBQ ����N�A�,0����r}��~UL�����/ZBi�6�9O(sJdJ�����C(�2�/L?��}v�<�����\�ku������糙O����	A|'��o�,e0>(tǮ�$�Zk���Q�_	j�|b�i��پH�</J����A(P���J_f�MW�f+��Oǔc;�����'���͑��z���k;[����!�tkG)/:�x��ČA��#��)�C�1��n��f3��_xET�G��b����K�c;n9��ފ��0ml��궁��O���hI���'�7�t͗��W��|��i�NI���D�DG�{��,�߄���LEu ��"y�w�"*��#Ux�
�^�03�����u�.��􉌣���Dz�^gb���V���ۻl���㏐�	�\X�����cv��������'xc�]f�]Bmɀ�6jо/��e'�)%B�VR���tg �x@�tc>�+��sT�<J��+N������D,$44A#�|�T��}�{s�ﺵ�I5�3�_��*A�XE��"y�%>>��-d���3��2=9��{����ۣ�\��'���umM]��Z�t)k���YvSt�oT�M���V�[{�,�b�K�m�f�0��Nhh�^�tz��l��M��~�Z^<S����={\�a�>m(�����w���prrbM_�`����oF��V���607c�!��{w����]?=u����<d��P�җב�"���v����}R���4�`c&J.`�WW+��};Kq9�x.��+�Eu��j6A]�vf������] �S\r�w�V��һ���Wa��>�@��Lm�C��]���F&���2�T�cl������s\V�����0dt,����Di6`gU�._6���\���Dp�M-ɩ���i��B744lu��nL\&i�B��IhvRB
��(G���47h\\S�JL߻�R��1��2_5���%��J`mzS�sK:3������ >�m�4���$��(t|�7��&��\��ac�؋n�v6�?�@y�A��'�tbNT����/y����bk��3�x[$��DȽ����a��x�_<�)_N��L� >��n���bџb�lY�,�/�����Z~p�����m]�;�F�]�}��D��fVb�'�8�]s��B꥓��땛�\{!�x=�Y�w!4�ch%�������N<���i�^�C���^����cIc#�נ��L�
�m;�P�\�8����GT\\L��F���v�ύ�\�W����\!D>�]O�:�`��~	��ϋ�3]���j����YD�K�������"����^��oE5�I0І���gU-�&��Dnv��M�7�X�2�ʳ�
5��U�%a�������rD���z3�^�����'&.��;��F���v��7wK;�&�����r�p����pjQ�-Ś 2��f1ck^չ�ݮԩ�p������a�r-or*$L~b��"������(eRh�g�`�C�p��.����o_���lh�#3� ���m�W>iî=t*a��A�
�ӁO�ɕQǺN�����En�I��bqR��O(�⧾��)�I��α����@��,��]��8vyT�w@�X�'H�!�2�w&'^B���F>��#|!
[�݅XW�bM�������v��cgO`IU��i���*,��w�Jg+@,0:g�T`,�#~8u�>�E��=�ѭS������Q���]r5�]�G����և	"���OUX���!��nz�4�`��Ru���	�J��ͬ��Je���h,K�xo��-~)�q̷H����KP�_�}���|��݀8����1=���+ۋX�D�f�vȧrj���*�>���&v��:4i���$m�W6� ^z�d�S�J�WD���B�5�-]���и5�e�k��\e%��e$L����}G�~;Y���R��ﴷh)
����/þY�P��T�rkޏ2Lg:D��.(�n��N�kBP_�w�ĒV��1"»����M��_�٩�����!Ƌ��
m������%�����������e��I�r�M���z��Y�qZ��}�������1�M0�m�]m�g�P��XS�g��}D��,�"H�:\#o9h��
$cvwwO�������D=�xa�����߃���};;��kR,�n����S/&`�=��~��"3nn|���hn`�m$�-��`�<a҂��|u�m�_4��p�y���=���gh���c�ϵ=��/�)m��b��B�6^Z\���]b��4ˆ[`����?������E�{} /5�(�dh�Z^0C]��J��6-�30�
C�����aX�w��y���`���$ۏ������+8Ecs�0iKAd)4n��y��Ҳ�@�#�����݅��B�'E��UI.Uы���wZ*�n�ak�Tj��J�V�'������&��4�7{ܐ2ZCο,%=��5��-��Ԯ%���V��g1�!�� F�� v�yl��FQ��q9JR~NX��Xo�]52q!����c��'6N�@o�{�.�k����w�530� uz��ї����K|�����Qٛ��4�#��^���}.N���at�4�ޜۓU�+�v||��E�i!������#*YD&�C��O4Z"�y�c�����,e�3���O�����d4g��p:��݆{�p;�Co��^~r���9�۞Ω��b���m_C��Ȏ'���>�.���Ѝ��I���������V"E=P����@+��Ũђ�L�0��`����KE&dbQ�2ƿ�g�3=H�vЎ6A��]�꭛�p�b�=��w��Lv9{M���Z$���o�������*���hn"G������%~�\���ӵ! �Ȏ>�8����M��| ��~#g؇���f[�YN]>$��!�M4r���.W|�z���f��^���3������d��o��m;[��l�Z�9������	�ttJ!t�:[��ۭ�blpuL[�4o����ɕ���L<#C���ۄї���s�<]���,+-!�			J�Ǔ�8�EZh�Z�,&LZPC�c�1�ɇG�34p4�;Y�畗�(Q��Ur���-^]�@�&,��*������jKY*���M\�8���;i9uvgr�1,k}����ԃU$�|�ڸ�9y���3�tȔ���������I��:��ɭ��n~�#c�@��_��fmM(���k�h�:�Y�Oo�?Hš��H�`�������6��0t�J��t?��{x����k�8J���7d��V���:;F��W�b�����ެH����XZ��ų��T.��FC2�!�nv���6 PE��)ۗkN�-�
w�u��H�4�0QB@@H)�mEY�+�[�ow��*(b�`��?�&B���.q��� ׻����QM`+�@�X�a-�V��d���Z�u|��[�P�5���mД�=�?���*�6W��\H�����~�5����@�_r.���p��FҢ��)<���lzX'	���57�ji��wi,�J�q��4���������]�ʽ?���?�:u�F1Vx�v�VY�.b�oL�շ�i�';l)!nQ���4�^o�"{b1�|�?���m���)@/��|��g��I5̗�W��G�&t�e�? Icf5�B�S#,��<��/�^4c�P��;� Wd��O�K�9璘�M:*Ǝ���o����H^x�Mp�)f,:>�'�G�ނ3�FF �Bt��9j���M�w����<bт�d��c�J
�^��|@�@�����:u{�dӎ���.�j�	�6�׌�֣E�}�}��n�\�;n0�ι3�i��e+آ'C�GҺi��XȒf!�G1�r�Q3��M��}
$���R��ȳ,J%Ô�&i�!�R!z9L�Bo<��B?Ԇ-r�,���d0�̃O�9<�
��	<\C���C'�����"�~V��Aztf���п�찤�tHou��(7��l=�A�|λ�XU[[X�i��.E�1tH/�[x,�1��������������Y�ڗS,�g��߷�Re8"#X 0�bi�E��o�fGS��4��W_�D�Q&�f|��e���i�2��Q��#���l�ᡉ�Yf^p��^=/E\
wYk�i�+����������侸sET7�>��J��,�v .B��G]-N�[=�;���ďf����OB[${�]������V���8у����� �3�輿�[{��cq��O�x��`F^��ۛ ���?RpId�F����)��ӄ/f�e�R�0�>�18ȹs����,�����
���¶@������_�����3)~���G����W4w�3�V3	�?�sܓ7�S�t�o�Z��~�!�_-�m�N��cW�nǑ��ܜ�O�Ժo�SO�� ���і�<����_Q!;@��6!=���ͣ=����#����^����U��L0��Q��Iܑ�\EHQے��� �sM�w(3�-��L.%^/p��'�%��A H%D��y��B�8�G�u�u3V�dj��V���S�9r�
�`a!��Y�n	_;Pz�v%��٪���*F��xR��MgX�i^����`|(��j� �Z�y�K=�� ���n�٘K��ć��e�a.�0F�\��6���蕋��)\uXP���"9Wz�.vu�U66,�	���>�.��|/������L�����6�����Ek'���kډ���%�#�C�:�j�LQ��zF��R{��eV�,)�i�x��'���"L�Bw3�6C&��t�ϒ��A\��"��;���v�غ`,�;��.k�]�H#Kge�뚥�<lo��d��>�;��ϛ���_�G�0�'l����=�q4{s�ب�<I�g��'�&��v�Gr�QAf�0�MGǾ뭱��q�m�w���>��^<) �[}>��
���u�YV�1uDt��#�z��Z���u�L�3�]�!Ru.�U�-�˹Gn�����SNj�ᠽ3,��G��Ȩ"c���^�8�0��.��z��Ơ�6r��!�B�c_�S{�qQz�'�}�N��9���cj&�X��-��i�L������-f��L�� �n[���Z~O7�Ʋ� �v���Un������������g��.'�V$�����5��K�q�	.UM�i��л?<uX��'V��\^�y��Bg%�Ã���<���0*oŔ�`��-O�o��\������~�5Ao�a�^�j��
>K�����K��	{��갨���ӹ����Hn����?��V5%0��#<Zl	��Ή��V��~6r�3��Sf��[�)m�M�8�����������kߩ�9��e׷����+�QB���
þ�]��@V!�7�$����Ha��9�B4��k�ۢU<<<~�W�P9vv�IC?��j�u�F͔��� ����T��v5	�&{d�U	
��fѻy��^	EC����%���*�SJ�,�S����s	p��;�!tΥ���A���=�O���"�]�7;��O.�����f��N ���|$����!�8gg��%L��Z��w=��=�uZ�0�b��pg�mF*�R.[W�8j�}Ey戵���v=�k��q��p�8j%��Їo!>���� ��V��eb��:����u�HQ����
-�iP�v^��^��+����0c���h!�D#��M|����OA3_��9��n�].�$r�FO��x��{��d'T��_9W�l�k�0g��ϵL)�sXu������B6O�� �p�EB�54�³E{6��GRb%�{0��M��w�W��7�%�	¨��Ò1�f^PpU�0��K��o���:e�n�?ݳH)r�̸^%���.�Z?~�5ۀ� JW~ܩG��T�|�xrr��Zvm��	V̏��� �'��&��:�^��O�3�Fi��z��1�U�d����ݏ����o��Yr�	x����N�h��@�ow�L�Y���xG�o���+�oڷ�p�!����)+YM�لZ�>#1��~0��=̽�:^�^��@Ƒ�L5��t�~��n�[dV�G��c �)|>�����'\��;�Et� �=�{��0�ݻ�`��]��'z�V�.'����Zi.}eS����H5�+�ɕ�:��� ���i�(����t����g	�����3(Y��x�&mUhS�CGdނ#��N�O�7߫b�Eo���UνB4��x�:�ÿ[ߗ� �_X@o�݉0�ie�q��� �%S��GtQrpZ	>1pn���_#���[�+�1�7���wu+̧�2�ߪv���f��x,�IB�>����X�K�l��$Y��
2�3�"�z�ڄ�2�&H.��('��W�4��%lp��h����t�V�������̓�{�,�b~~�Ɍ�֪����~̀��yS
>�L"�r��)�}�B3��bC���/����qm�>�o��d�wᮽ�t�u_���#�3���{4~�����G�%m��)Z���D��.�1�s5J�c��]jg�L�����H'Ӛz����(��&�����lL���A!�F7��I�Gzzp^��KN��^Ճ�b����S�b9��l���&-�NWs�x'c:����Q���v ����\4��S&�1�su��]�.]�/�C�j����Ą�@k����@�c����#�+';���9>y��¶�ٜ��jPoÙ5:Kz���gڕ���c��{f4����C��LU��MM]��LE�O{▛Z��v�տ���Ψ��L��@�K�'4S!����h��W���:��VRG0��k�b�<%����O�Wkjj
��6*!g��7/�f�lJ�7N�񎼌O妹�K2&�0���*������"y�d�����J5Z`'�,F�--�~�"���_���� ݑ�ʍ���b��Gw�&����W?g��G�+]sg|o������2Y��Faݜ�V;g�t�0�D���<��hg:�S-1Y<�Y��c��$������ݲ�����ɣ�d�n���g6�7g��I��~Y��:O8�GPs���ǥ{��a`�擊q-X98��vJ�HCa��.�y�1�5��b#O�匙>��AL�m#�ֈ��8�8΍�s2c�����S��J �a�n��Հ��q��cC�n�4:ꞟZ��Qݼ���ڹ�e��3�"��q���g����e��x7F����-�7��*�ޙmVn/�M�MvЏ�7Jvu[�p���>äiP10�Um�ژ�4	�n=:����P��Z`/�D����_ ,p��r�q��l���W�10�gg��2d�z�|!��3�as�E��d�����r|||]��V&zM���ۿ)Q��ey.��������g�[)�X���sU�o=.)����cJ~���m���L-&����B��Ń�H��v�M\���<�_1�7|[��ɵ�=
'!���!��(o��ރ���X��o2
��Ռ�S��r�\N:^�Μ���/)��%a�� �|*�<z����#Y"�YZ���J� ���^�;�F���>Oΰ�mgH�4ML:�d�?���d��Ì��-kS�J�t�Ċ(p윝�|�	�Srk��>a�n�4��X��S����qdV<D)6(V+��C�3]���^���+dJ��J��ޅҷ_���ג2m�V�b�[�%0���1c=Η�igAf+b	���N��?�-��J�<�;F#�k�N�Z������5�	�ق��6y�~3�JXp�z�ݑ}�L��d�y�a���H��=��E���ۋ.*�����~G��)+-����~{�7���G����=y��E,&�VX�6<���[h�)Y�nts��m5k�"�h_ؽJ�������51��	w2F��{$�G���t�[���zэ:����qK���i�:��/J�j1�ªƓ9��K�g)tp�{�<.����y�T���H�'x���1z�=�	1���^����V�oJ/Q�����F��rU���ɚS�ݿ�t�t�S��(gl\l�+H������su_����m�m�c��j2��+�=�YM�^��������g/t��Y�Yپ�}{�U)t�<mngٟ�	*?�$����kb����,}䨠q۷"4zd��4~��g��yzT�b�
�%,՟e��C�l麋��h�W30h������g�jB� ^]ڏ,�5��kc@+�f���S�"������cMZ�ىv�&�ޤ������[ۖq����CZB���iiDD�AJ��A��S��:�O<��?���{���/�.�����Ŏ�د�/ɞ���h�D����ǹM��?v>��F0��Q�pAt�5��s+�c�� �_p�G�,�5L���p�P�*Grn�Y�;S��E�q��|��bI|@�c���2o�]��g,�MF��=u�ae���0-(�L�����^A��̹�����T�'tT��j�)����wciY�H)<A�&�3�� �Y$;Isp��)�ؾ���fۭ��W�c[[[�F%-����_Zz���B}o�Ů"w�����M{3^���	]�Ѯws���n1'�
��t&��Bv��*������c��}�\=�6��,�9�{,Lsϓ*�g���-��{)|�D��|1M'�S�pA��N��$$�	�l�^g,����]�E�ڸ���%�4��gO�oT���+����w3W�s�A�G"UN)��t|S�"���õe��
#?L�'0���u�[[������IHHpv7�#\�C_��Є'���G��q�r������,�sC��3tց0�7{����3��"]����,���%2�'A��X��������	��A���;��f/��Wލ�cR�nA�B�j�t�V9RU��d8� @u���;{2�7���7A�'��*��@'�#��T:�8����G�iq$.6ؿHC`Ⱥ�p��Zپ�K�Z�0ޞd(��4��A�/L�D4��R�9r�jBLHP����0˙��uPؖ��vן�e�=4�ϣ��.K�M���}h�a�W�[��6����U����Պ�N��#8�)�G�����Gz�D��a\���jii��1�cO�1R�E�_�� ���|~�������T)#�K���x���=9<T�r=���_)O�僷�	�����	#��6+�q�L�"@HT���Sh�Z��$N��;w�#]]�n���t�Ⴖ����ʡ�F���C�	���7-Cx<{7��m.���|ŭ|O><�Oy�r�)oY�Q>o#N�4��+A˾�j}?HbЙ��>����9�_���=f��5bE��3���O�����te�����_6�\X-��NNN�oK:���Չ��,��s*�"�
Њ��0Z	q�#g�
��"(}������$"��2�ں:¨�)�c�HT�!%�+l�ř��jLV�		��;(���=v$)�e��#��x��������@Z������+Ŵ����҇LE����~㟌Agm����4�%$�i¹]�����ņ�>��~1��ڠ(�O�9�.$f�V^o�i1<K������3�}M��IU^/�Wof+v�t�F�TMG­�7��-�P�"�QO��앋��Α�a���/Y4I"���h��P�)w�n�u������d�l)�V[�#qUzh�e����f�� �|����ȜW�1��z4�_;��c��E.��	G��.)b����6�,��( dg23B�6�w�A�O�&�r�)�W]�A�Dr;)G)|����~T@< ���x��-ʁ��R�`[�6�D������vA��Kղ��e�hs/D�	n�.nh|�l��A��L��\��Xf�軞(t���&�S��n��jH�;.YMg�vرo]�ni27�/��i�
ߞ�T���3���)k�y0��)�����}��������B;�w�'h���6J>~�&�I���������`WD�Lx�,�V�;�D���sRR�tK&\�q0\n��S.|N��/s"���R<�1���W19)������t�߾&!�%��̬i��U(r��(�y:�M9m�6v��v���h���
n(�50��),��r��]@�/����8��z�g��4���J��zg�/�7���P��(�W)�P��J~�8w6��xFD��3ì����ڠT!^�GI�˸��['a�4�mo�J%!nQ'm���yo��Z��_/9� �t��N�%M�%	*9�V~�p�>ɟ�`�	7����4
p|ټ|�xgK��3�ʹ����W���a���!��m}}=�r{^�X��-�����R.��ke�`j��z�l�'="������u�z�_~JG��i�W���<�f��pC���.��%�[�^t����A��l�?-��������J������nư�ȑtط�������n�������?���>(Fo��ܨ�f�+l��ݍ��Γ�)	�ٶ-D�ow�6|O����W��w����;�6<'�YT�q�/Y)��i0�	�ݘ���tb���WE��'ߦ/����;y����6Iľz���#i�Wp��08��8�U\,��^���+��.���K��>"�w4���%e8}���{d��X�a7���`�{NG���0�h]��h�Z` >	|yW���e��U���q7c`&Y�Ǐ{>=�����*e(�߿�x�_�����������}-y��]BY_�-5�!,���U(\+��meF��ťV�X���<��ddn�%�M9.���O�5��'�Z:B�0�~	i����b*�E^�)��o�H��CJ�k�3�_�Yi�c@8%�1�Y�g����b�e��M|I�1C��l�К��=oɁ┇���>��eB����*���'D�y>ʀSix��y�
��'Z��ѼN#'�W��u��eQ�Aԅ�G+��ʷ�o�;-^��	jB��~I����Qk�TTX�Y��h�d�����9�g��3Y4񬬑�&x��;�;$R:~��"<�����~ٴ��gI�:+F����d�lkml<����>��i����^��q�8r��m�h�g+e�Yąa��(9��C��$M�n���TY�.�qi.@��6���Z2�ٹzl���W@����-������ࠦ i)�W 6��_U�st�[)n�n��su h�O��w�
���+�*�Y�<ěE(�/�\K�2@Q%��D%�����~��eQ1�$r�G�M6٠��M[[�x���\��e[��UH�Ae#���u3���� aP��Ǒ��i�{}��3���ق��P���P��O�C΂�Yh��K���j� T\����S<&�g�g@jEӮ����^�P�crYH�-`cҷ�ˆm��l]r���D�9�^�*CL&Q�s����b�����$Z7r��^^��ݥ�cc�������P��BՖ�����o��o�����ʑ'
5������,E!�����Xn<7
�|��eJ�ۄ'5���\@Q�na�Fb!ҳ�
Nk���K-�E�r6�N���T�n��/
\���O�ؘyJ/֎'�����!���~xx(�6�0?��o=ȵw:��G��w�p�ŀܰ����K��	������++�3�~�3�fvRJ�ţ���D�H���Hp��%/��)��9�D�}�E:�ā���M����fe���I�&bO�:�?0ax4��A6F�%���[��v�u.�)AС�����Q�MÉb|ċ��n�����Lm`?@
h��^�^Mf8�3�B��LFrQ`)|���<��`�ɝ��iT�|wkKI�j}�vZ�Q��P���4I���������)�j�����G�T$oE�ZG$�6��ʻ�iPꊌⵉ��X�$��@8���n�D9	K-ɸե��;����)TTn�C�*��@��q��*mm�8{��`q�j����S�2=ݗ��x} �/Jሯ���r��o5[�W}��ms{� �T���t����c�At1�uD��(PiTB	{ܖ�xA�����[�5���j��L���x�w^�6��4�pN��Kl�,�v2��>����r
�[�p�m�(�Y��g�X���7�gEi��9J�4��E�"��.��6�1nq�	I/
7T|���s	�^�Ъϱ�>�ܕ�GX R�4���p@o�����F���*�f�#��5,mT.}�)�*��g�\��p`�>�D���˫����{F
�� �Ǵ�U¹�:�$��ٍP�������:�y��ŵD��YHQWmBe#j޾In�H�|8��ðZ�+*��C�#ѻ���j~��۠��ǣ�U[_��Tk�م�
�T��kL�p�Y���M.���,y�k�,�D�n��<0 ��C{i*����G0�i��I�Xx���3��P������?������אq6�[�K*�x�sjxJX��"� ����<�O8l�H�<�ؿ���23��q����|NM�w
ц/��_���:E���P��@T���af�b��b����U.T}��JM	�J�p5�.T���~�ө<��H����4�' �m���k��k�M�}_��OÇ��:�oF���I}i�`���� ׃��N���4`���!6',}����]]�|�<V~���3` �Xݍ�ꂶi~�����tS�ˣ�	�ѳ��wM�F:>��o�"��$Sv+��͟f��&
�5�o���'*_ǲ��К��/�y�����O��4�)TF$_�񭱊���¸�����I�P�#Έu����_�GͪK��T��A<��.�p���\WS۾<��H�`CKF��Vg�>Q�y?�c�T��ķ?��tmW:�6�(8;���;�mxG��)z�����ㇱN>۾�B���m�B�㼘���Q��N��6ڐn�w�N�f�ۭ�l=5s�8�T��޷��͍���f�4G�]�~�A^�:���88|U�X��K���' 鯛4m�����f��5y,�^���՞��������V���Q�����������<�+�	��^l_����<f�L����s��HD`�Xl���.NNSW��F�����K.�]l-����Lx��
)��[C�Cr���>Ɍ��yC�蛝}�dDV��x�|��N��=Pa�l#��V�2=���Ϗ�^�C<�,��u̕�瑗����_��Ēr�R�?U��[Üihi�#/���4u��;���\?���bb��ɲ�}���t��k��}������'��{3FlN�s/��_��K�:�'�}�y�#^I�e��R㍝��#�Y4.�E	��]n%HN��t�=�L���!Z�d��Ί� X�Fl��W�K����6��8���R@ \�X��K<�����nPD�@�z��H�Y��ڥ-�{���t�E���ߌ�g�<!Y���r�E�&���@ iCp�'�eyGy%����E���7��E��� ������~��0�^��PD��Z��%j�{X�.⤈��v�T�8����=��ĳus�<�����^�P���!�Q;���<;2\����1���ž&��dH�Z϶l������7���ȟ�}��o�˘8T�|���$"z{]�0�7R댉=��E���[ϳ��}����b�P�S:����T���N*��+9xg�۶�V�x�k=97�w,Ufp*Õ�J���;�3��\x4:`�G��P�?��Iڠ�M&nW�z�v���1�hkl��_b؋�~��*M㎨	�W/��S����«~���m���b8���~\Q���G�K
����9�1ڔ�%z�Wg��W~X��`����V��{���hmJI�����A��]O�R��o�-���B=���`��(��CM�<�@f��ej�������^�0^��0���.V�Z���u�c+�$7R�p���w��V��եQ�<�츁P]or���׿Z)�R�{o��Y���t�oI)��-����3S�S�WD6�0�~ݢ���������Luy����T��3��G@�9@��#��~Ijћٵ�AI�(����.�-����Ǐ��7"�����o�[�x����'s���:�������XkeHSh9M��}�y�:���ȪZv��W�u���w�6#mӃ�m����l(�CߵvΔS���Yi�GՏ"�c3��^(W_ή쫡��HL^��\I$����aĄ��@����wę����v���<"��Aɍ$���qPoI�ڧf��ͫ�=<<��o�~&�鯑��$-�U��w�%\]�o���&�3������F~���~
�A����u�����U�s��x��}���#@��(6HU���Wz��W��bKf�@��5�>\,�l�vO�ψ���qTh���vw"���5��	6�7�/c����q���L�ߥ�$����1>�ԫk|n�KU���"��9�}���拥v�'��aǁ�ȿ	���Q�0B�>VAL��(�1�?�c��l�`�(De�ܣ���7oG���X'h?}3���S�զK/�$��	tWrف%��A"���'.=�2ŹF��4�u��(Q=�^�q��Y��=Ԅ]���YY�x�L��S��1}yY��#ĦJ���:��Ҫ�g�/�6�r�k��"�*{-�?p�wS�p%!kZ4����%%�?ږ&���DA��c~S'����P� }���r�D�N�Ƽu*Ґ+-�������^�b�<�Sa��\����"��E�(�F,$3O4xIHs�9��ʦ'�e㧅�t��q}���c�J���?υ+U���0_Ɵ?Ǣ����Z9���+��6�Lz�	R��� �9��� �n7��.�U|��|�Mԥ[�N�����a�_*X��x�L��Vo��n�d����ҞxN���] ߆��.��;Qj�E���������#�G���=�垈�}D�bP��҉�=�t�rB�Ɩ�rDx<t77E�o&�m�5
=��3 ��/d .��BN�����������s/8t���ܗ�	:�����7�n�Z�l|�|����x.��~cc*�7�G��t�e����Iǹ�R�U, �) ���$�����cߘ����Da��V�L���ؠ+O]��N]x��AJUY/	�.�U�闼J��`��&�x`��g�L���t׆���2,o�`)f1�t&Mh�{{��9x1Y�8��i����+�J��	�M4��GR<����Cg	M��e�.S�}ֳ!e��8>>���X����v��w�1��gS�:H��BR���qQA���#,��U�|�*�᩹an�jl3��R9YW�e\��(�������e�Ĺ�D��D������|ё�3N.�<����W8��!4��8�j�@被O���0n���l5-���r vu/j�$M�@$&?�G���y����fJ��(#����v��t�ŏb����=���L�QD
�l�12M��|���Zr��|���>��3�'�Ҩq�2��<�p@ܳ�)ډ� �~t�_���P �Y�����(VD����n䠳��`q�R{���e�n�Jkbr.��2}���(w�@ ("��V�hh�zq� ����z<�y�Z���(�3@�����8j(�n%7����,�IXa�r�/p��`{���B��,�'����\�ʳ{�� �u �P� ���^�^x畱�R�=��Vj�Mju+[�:N,���!��!^�!4ש��GO�nX��9�%�b��ͫ�0!��m�'�b�TS�Y�k5.�6�m<�a-�,�k�D 5�/�H�4JZZ%~8�׉pܿ�J�6ZC�Ё.�U#�����'��Oڶ��z��a��z?��Y
��$N X'��¯�#��)�U(�7Ӓ�;��3
�3M�AԺ�� ���P�	�p[����n�r��*��&F>��:���	��F"M�h����\N!�����"����)�8_D�&�~k�h�t�L/��	1n߂��js�R�ς\k�e8�8�Hd
Z��_��u=V
��Ąs@�m�_떻M�j\�lTt�"hR��ۼ`�V����kl2<�SY�_:�����v�F����KX�o�%�+�ϛ�{?��;XU�\��ö	l��b�&YQ�%'J��TM��)+�w��G�*C��<5�"{L*+\D���~�-�s�֒ߖ.=Sʨ��Qd�(Z4�L"L^zA�K�ԅyQ�����6�?���2p���r��g'4���2Ew�<���±�(��y�h�VW�����'�):\���?�湯%^��O�iŲ��
�dEǷu����m�PL���C1�/�����t�6>�9�N���難G�5���@(6�����yYT,Mc�=;7Wt��J��O��$;T�rI0U=?u�v����{��k�n俕�/��?�:OL��@�p��H�,ҙ[Gɦ�]״�������=}�-9�!���w��5
�\=�\��>^�o1��6����/
�__��R�">�T��RU��yb�qMcZ�~WuӼ�m�i�8.�қyJ��qt��%;�;L{�эFCiڦP�MN�q�y�����mK�,쭭�>!W��bg��B�!]_n��ػ�q+�.Ur(Ce����sGmcR�����O��ќ����.Ι��{㞏��}�e�V��C����㗯zP.s�9v��xX��(���\���[�-����N@� ��)'K�P����m��r��އة��m���n���\����KH�BH�:zgE��_:p�������D�K�A���+�L�ѕ\�:����#����@<�"�G�(Ж�'�X���ī�덱~�g:qp�,%-����wt�ms�^�,�d8G	�Dg�V7ߧ0�qԐ�ܔ�Q��ل�8>ߒIN��)�SUU�6�.��*�������e�H�����XO��$���HP ��!m���mJ�Zc!7P;3 ٻ��F%�pS��~������� �ɤƾ`צVS���O%�P�!�-t��M�8ҖW��R�U��I�dJ^c�M�V�n*���k"O�C�����l"`�}]Bc����\�'T�ꬍ���`#�'{���y��U3�����^���?%��E�l壖bI�ƿ��\��	�H�:���ӿ]�0�#������F�����储��y�`'ح�f���u����
3�
 ��Vna��Ǉ��į
2pb�x��XS�V��m�$*����k�a)J6�U��=�ӂ�^/^�*ZJ4G��8j�;��[�*%ԇ0�~��c�0�~���y�<���]|�:i۫zX[_O����_�-���*�Q)<���uϕ���z�\��*[��mZ�!(�a<�n��NG�K�v��d��I���a!O"Z�{�� �]t�"s�S*]��\�͂��G�'+Xܨ]9�m}b�E���L�8��0I��ի�sy2n`�[���d�R,�O{ۿ�,
P�0���<��I�4OX�fN$E��MH���lK�Ol����+�kaQަlT]D��B�)����� ��3g���Y^�����F��8����</ܞ�W�Ws�R|���_=sO�J�$�9��ໂ�!���q���X#w���3��QT��zҘuj�l�A-^u�wRu\�����e���R��ޫM��M�-�M������3�^�p�<	M�߼���Z�V�0��� >����%J��?}I�m��9+L���3�s�A:��!�,V�����-�a��8����u�1�Z&����w�xVUwo�w��e��@d�r��=�nV�k�\���ɩ���7�M�yi�>�6�.C�>�U���渨)�bT *���}�����ːhR2��nI@	X���l�lm��)T=�sS�o;9y;@�)�������=y�AJz�Y�K9w_P�׽咸+uB�� xxx��{��޶�k���5�h�'�Ny!^�Q���!��.Ka���N�����>~O��l��(��ϯ#!Y�L�c���Of�Ԕmll�f}��e-hq0�z���**�|��:��owI+�h]R�HH���}���{8}yZ���JO���}�:S7T�^k-��f��HK��֢j�v�V�� �`q�j>ĥHjuiiإBX�!���N��V���u\Y&�B��
w�o{��z ��0H���(�g�r�w�ծ_��u��<'W17?�s���-'�<<266;%��y�#H�+�ۼ+��u怎���`Wv���I�](�
d粝k$�a�~ �Ԋ[�o�n3��CHo/w���vڬ���ϴ�A`i��G�����F�� 	�'HZ�WڗQ���?=Ȟb`�f�eb�Q=�U�s�q&bj �����*TqCgu�Me+�>���
[�i����`��'Ml���ɨ�U#w�����\�q�.�j�>�ڡ�Y�7���R�$��\�>�b'P��))��ev���%N$��Q�
�.}�_B��y�6��䌝B�J�j��v��/+9�E�Vma��;���)�xm��>0�<Z��3W��3�����K���AEX�Eg֘�b�9⻩�����y/��M�}�볲(ʛPL�fm�k��=�ӏ�=[G<����f$0
�V�e< ���[y�	ҵ�� D �]P��P }	�ߚ�ٽUR�(�X�kc�\�F��a�?�20x�q1�ͯ�LS�jf���8��19��/{n�g�da��vi�<\)����c����te���o�3k{=�V��鳬�ݙ_�I��*oOOOO9u��|gl;�6�}5E����=��|�'X�.g=ex�y� ���C4Y �����*����QX,wf�g3��^��q�����
0�h1�d\���:
�m����.YD��V9�U��/�Z�®H�f��B���St!.9]��!���$���]��?e|MO��MsZ�i�,1����X�;�Q��eʞ\��3�0'̦mD'ШL�m��2���G��-5w�̩W{C������y>t`|=n�:Jc����,#�X^>!j�[�~F����� ��%��tq+R��	�N�m7eLk�oǬ����K{?E��v>&���4b$�f�2$N-�)��ɵ>�� ⟙�(Kjw���+��w�������uU�����1ǖ���$�EGIU��aǂ����0F�B������x��GWQ�{ �[�7A��eg���T�1�Җx;�{���
OT~���)��0ǫ������ch�-D�?[G���o��ӉaMY�� ;:ęy�Z~Y)��u댿�
��8nF�K�rvd%�E]�fͬ�XL�*B.p��!��p_|�o�re�0Ȣɴv�C'ٌ9�b(!aJË�jgeBf �#)�8Jl'�򩩩����;�=�TtAi���V��0�Z�L���ŝ���Mdqd�ko
y��?�����N��Ts)2���,V?�?� ��u�>���P�C�v�Adu8B	�r�b���3-y�����*|#�Z�s� �D S��ue���2]�]�4�\]B�5<��!��א���(�Ly&�ز��LE.�����cQC8^́��t���q�c�1guMk�^d��5	��xQ]�uK+��w�����ƈu{�@�X���lʭ���5LDv:T����cޖ ���^����]'�i�c2��� 5H� �urҨ���;s��]��]����eQ�E$��S�F��N�E������%m�>&�p�B���Or	��gg�C�(+� �e�9����m�x����QҢ�`����b�Ω3�C�I�?���k����]_����T�;�ҏ5�ԥ���y���K�X������׌�{�Ɨ����&d"d	����Z�ꋃ�eOo��B�X�)Y7�[���l��+����@Y�@����$�m|��?I���T���O�$��(U�<q�u�j�/-��$Ҭ�)�R�z#ZЬR0)޻C��%<z�#�}O�#���c���4�8�n�y��&�j�n� Z����^�ƿ���,Y�L�+�(���N���&p4C�Ԇ�a���&��L�صd���w�F�r��Avd7Զ���,�L�o9@;������4�2�����y�4�Ԛ�%}l�OÛ�v9,Ӭ��r�3c�����O���Z&�@��P�Dx��I�E���G�~H��+����kwɻ	aa)�8@w����~/N^�tp��njx��6n�
rA�>���L���v����Am�b�_�æu�r���Q�h��3N��A@��m�9}�<s7���㵳���={���Bh�y9�_i�d�����*瓏p����5�/-^SAY_,L���D]ˠ?�l�����N]	R�W=P���t�g�������[>�1�o8�\z�E����'ކ��53��!%[A�n�*�9��}��;u�iD��^Rfxn#T�Y���#�^c+�Zq��1[K#��y���fim� G��,A욆I��>Sva���]r��o*?,�d�Ǎ;�9���X"�ơv���U/�����D�C]���f~"��ӆmg;D���[ޫ5ﻗ���Z4����j�k4�}{5������r�����v�|��آe�t�{�\��3P�|@˹��Uʎ�FY���"*\�g���RQ]�L�!B����'�y�UNn΋�݅;o�@Ѯ���6��J�@Yb��QD���	uu�$$�f���a�9��W�^��)ޮ�	�A4~�>]r�uPz�?���4�0[~�E�uzg�f�E������m�揽���z�1���V25@�H�6�T�厂;"n����=
H�O�W>�l���w	4N���-r��p��wz8Ih�8�އ5�a�|��٫�bv��M*��-�c�i�*�S����	D��!����N+���`�/�$@�1�U_�L9+���q�kg�'��6�������m^��TJ(��Al��8��|K�O%��L*`���Z�ˣ�x|���c6���Ӱ��o�e趤�~����� �������V����x,��NN��w�� ?
FM�[���1�����P����)#rH�O@���)�J�cخTlm�:*��F���z�G^X�W<_�z�]v;ċgY"iL�O�j�>�������p���qw���\�w�{�X���ȝ&H=���lJ�j��T�x��i�L4�QZ�\^_�C>��f$Tn�u];k�_���}*���RM�/��s^�O}`ތ9�^J&�8��{�:S6,�㑨�\�@]R)�B�s���l�ϳ_���zn�o�������Ev8C@g𾭧F0�����JsUF�9Vw�O}9M$#|ww�"�T;uJĩ���O1N�
C<u*��Wѧ��FJG'5���u������M*3����8��|J9R� ��R���h�M=�����::��U!%��o�`�
`x0���x]:2�
;�<Ps��o���[T�[��r�9]7�k/%�sj[�Z=���/m�
�v�"�Y����0z¯c[t�
��^o�L
Uw*@�ؗ�N޻�:�@(]�1f��뮵z�P1e��?���q �06>�j���B����;N/-��]�7��[Q�	���N����/���KYF"���k��=9�l�$�K��@lj/?��m��$`��)��о�<�b8v��f��v1}
�['����c�R�G��X�P�N\�t��������J?\� ��p��Z��1t�:���#��ީ����fu���� ���0783��C��i3o#����nC�ӂU���o\�t�Q�ߗ%�#�&a��vc|�[N��FQ����w�:��x��ׇR�#0�^�P�l��DʨN� u�f�y�!�x�+�WX��e��)�DTڅ�����on�6��.|ե�"�B��S�cDr]z�c������4��r���
co	>���H�+E�Z/��������Ȫ���**T_H��#��y�T�]h\өH�q0`ĩ2�εi�����T�6�xp�i��J$�?`������'b�{A§>sHU��R{�iӛ���j)�f�޳����s�oy;�Nz�q�M6�Ki�36�4�6ʮzŋ[Y/�����i�����g>.�p�@G�劖�]�*@�ɇ�G�9�b��02x�:������a�I;�rN��ɘ[�>��3�HXJ��N�t��k;}���͐��$�S(v�~>?���k:cN,��3���h�"���hbWC�:�y���7߾3�M�7�T��=]�>O��;�O�5W }��%g((E⺭[�U�
������o����^(+��tG�;�����~����B���O`x�4u��%7W|c0yU΢���'od�[oԨ%�1�ʱ��b�o��1������O�'r߲ؤ�k�=Pf��p#�.x�6�4^��Dķ*n�0�!���E*�~-��ޛˎ?rA?���k&�9�HNv�?�BGr�٦,6�'Q� <-қ�B(#!L���~�m�"^)�ޣ��j�"��T�;����J�̆�����4s��D�ƈӉ��q*׺L����e�_ ����HNќ��y/�&N2�j�6��Q���E��4xΧU��3�w�$�	~���Y����K����{L]���4�|���Qb�.��[�`��6a6\�dﾫ�~��y�����i���.��j
��8>6k�g���KX�F���9T��&8�8�����{{{�ȫ���5%��g��� ��rs�.҈[yb�^.�L0�ܤQㆅL�L�̎{�B�|��_�S�c�ȭ�*Vu~��-��6
;v�4j��ˁ����`��}�����/��O
FCgo[��H��_��g��3y���y��&Sp�Auc����ψt�>p�9""����:�]�8Kz���`�r���s�ӎLLP�����0	�nI�t�سmm��g���U#K˂�o�u������W�>ڼb�95+�H�h�����̕��߃�>Ɍ�2ݶU���jP�v|ƾ�&����l���"���&�!��u���Џo�{�8���<��ޚ�Z������iUm��%"�0DZc8J��%z{L��A)�%X�u��c��G>�(c,�#�t����wMh#��H���]g~����3{*�s�@�oedkk�)�J�+��ч篼vʄ:�t�,r***�p����R�L�;�X�z�kL�q��X�d��x��6�" cP.JH��<����፝*�b�.2_�k��
�M�7�Q���-��26��b�+���|8�o�:%�xw%Ƴ�Mq[w!d�`On8�Rf �ч����f3�����"�/`C-ʦ�ԭ��շ�CӬ��ꧮ��獘7u��xzNFQ���b�p�la��x�6�ͦ6�.'�����{�i�Us㍵G`�r�I����Q?o�w��AȘ`�����㦵�(���Y���w�A���5`@Njpz�3�� 	dc�1�^'U$	l����%��F�ޤ_yl�K�w�6]�V���{�'��ּOn]�(`f���϶��i�0|:�p�+U����&�ѽ� �W4m�J9�1BU{B�#�7��F��a8��cO�=%���l�q�c��0!� �>���*��XD�T]�4��N�zK�����ڣu�І�Iz�������\�~�q�h�wX�&����ss�_��7�_��Жš��	�$��z��{���d�������"ls�H	���Ȗs���@AF��cI�'ᘮ��B�Ѭ�xj�Em��>Bךoe��0
*�˰o\�����I��1�������M���a�=uE��",��r��E��A���˄?*���E�D>�?�>c݊�s\@ix`�5�G��K��5]7�B�`��δ��v�t-5�!^W�b�#�]�4�&ح7���N�eW�2K����(���8�@�<Yp��; 9�lXHO�@Mǀz&���j=�t�a��[��5��b��C�$U�svfC�XbOB^���<��4�y4Kd������}�p�//L��7��?��4�����ʾQ<����{i�z�P�3�t��L��c����)��_�`9�#?�[t��%�)��) ���/{2����I�i ���P�v`g��O��X|"%�'�g<X�g(l��J��6︬�Z���?��E�,���ð�*��'��fK'���+��s����C���%���N��h�]�r\�[i�t�+�R߸�+ ���9��;n\!���X�6�"�@�~�us��&ŢqlDs�p�Kj����m;Ϲ��o���Or�0|+:��I[��!��vt�<8�@��UB�T�G	A�A+`�^� ���,L|bbU"U��	�-́���/o��DVR�+�r��l��$]*�\�~�̗�ݖ���ܰ�#hhud��F��Oko�l���y�tߏ�2�BXS��o���J��z �qf^6��m{��$e��d�
���5�=�%{����x�~�2��U��g-3q~P�<�\ay�u��vf0y��oNj�e��fTV��>����+,���=Md�#	�E�z�@���B���$�Az�����'�#��p��&r�M��߱��k�������nʗvRRN�C��D��&K1d.�@���r)���,��f�*��࡞#݉l���@�oO��v~�����l��S/]�@����j F����u��z�u��\�b`��)*4z�o&�"��?"�"ֈ>%D�n�pp;�	l���-}��_fr���&E�EP4,�d��}V��xz�����Y����.���C���]-2+��\�a�ծ�m�ej= z�)���@���@�fb�R3�dmwW�6U�u�T_�
U�����KK,ͬ��ZY$��K�rQ��m�ڱ�5U6d1�U�������1�*�P;�`�K���r�]�0l�����!1�L��>�s��.b���K\[���`_�N�~T���#"����!��r�g��z�?��6��TT��3�gޔ �p�w��_A��$?������L�5��S�f��؇|	
N�}�^�5����]���ӆ�q�L������P;��1i��n��~U_B�~���'�Ly���ӭ�����}�����l�\C�'�7]��
���/EX�S��E��|sPF��]���?Ŋ�$8$#t"�)[ۺ�_�`i���{�\]����`P�7©('n���.�ck:�6"�Y=*��<�pRą%+��ҟ�c�_���榁��C7+E�QfH�+��{��L�C�Q��;�ȍ!Sv��+)Q
���)��P��$h�%3��-�_;�����G %��X���6%}�S������C�\H����%$sӶm:�S��|9 ���kʍ���(�:��L��)�[�8�X׍M'�d��z�Zʶ�ۤ��f�%��}�K�-�-�?ItKd�������k�:�}����3^��']�a�-^�qf���鯪�ϝ�._.�%;�t������9]��_�mj�\�w��}uXT_׶���� !-�"!ҥ�! �� ݡJ�t*��-�1tÀt004|g|���^����ǹfgf�Y{�{�k��q\������ �T���܌���z���/����{�+�O���/|%�\[�-�|���T�	p�>�A������*��f����;(a�n{���,*�#]� KN��ˤc�,�'�yg ��)ѱwM����xXLz�G��u�ꝕ3E����3N�)5���������q��˗3��n� >�Ƚ&.�\t{�	�_�%��{h�r���n˹�m�:}� �}�࠳@�F�c1�ss!�};B���9s��u���C���d+A%����Y\�6Qf5����JK�>hß����ق%���?K�氁�d���viA�@F=��I��az�qTgpC%N������Nǋ�cyq\�q8�ZS�ϴ^?L�MM��Ծ�=(��NU;97K�JXI��w�I�J������*s�49��S���-I�)��NC� D��CI���0A��T�Ь��H����g6��{���t�}�ٴ�*�^����8��c��\2�z
���U�۟i���2�Y5���8ǐ��������0�O�8��L�`�yUn1�u[`�஫�ͦ5�󓃽O	���if19yL)X@crr��o�}�ҫ?�h�1A��M9p����i��%G'��@ Pa1g�qK�`c�Ɓ{ǰ����]�=���z�dC"C�y�������U���1�o����f��E����N�d�W,H��)��>� ��ټ����>��������єV�/��&�'W<9If[!�pEo��RBP�{.��P�x>z��K�7���[=�ho]-�5��gX�`E��?� ){nj�N���EG
Д2����'�5�pJ�˽L�|'P�h��F���8w͛������l��
V�%LLV�j޸?G!��V+1���S_ ��7��7�����5��r��W�e�#�oދ�.�3�ȭ�&QN{�{`3CCk���4�T4CkS������^,�?�_���\M��[qxG��3e���w�|�$��Z�@Ժ�5gS�tK�5���Kآ`���b�3Ȣ�wѤ�"���@,vܮxL{r�d���I�kй��0�S
`��"�~��˕�~&�X!_U:�NS�k��|I��6���^�.m�nS��CF;_n4�����e�
2i�To��Bj@nݜ(mj�9�,�X*M=��q����T��f9Y&�X#��]�&��ŵ�Tr���/���y'%���M�-MF��=�Τ!����Md	�i[' 1h��g���x��������P�S�D���h<�[Txz_�^'���z^��.]x9	Ao�k�hc��P^n|�HMr��a �ٻ�D����6�Gv4�Y��o���"
��d��|�v(�)�T�j4o�iL�j_�Z�m�� e�2	������;�V�M���N����/U�����?���Tea�r���h�]'Mla��3++Ǌ7�I�M�n��� 4�[RM�8�äTTbݴ*��G�e?R�|K��|��Y!��W:mo��������fq|�_����e(t�I$e�����8�mcA� x
~7���Jo�������.�
f�T��	F
����.Ȭ���@:��>$״�G>@�H;u~��+����NFW\/�Dɋ�ܗ]��.�}G���j�Ѹ�C�˙�ۃ��^��k6�kF{�,Q��~�n�'���I���7u�m��I��ؿ������2uщC*�z�1�}OE�*�l�.k:���Ζ���Ҕ��`y$+�K���gffo����*��[���?�%\��{��.���E^�4������n�rzi��p��
N�S0H���1���¿�eۛ�ֻ�M6��{&�Nߖ�l��Yq;�+��_VtD�s��qi�3hi��lR�^�'bi�vm-�o��>�^�c�����%^\��t�"y��C))���ɲ��'	K��:�#r�����&S�f��ں�n/�ڤ3��ۯ����ď�n/J@�~ߦ=���x	��j�{BP�dk�u��J_��)��Ykཽ������J^��;��7��(�N�mn�Rr2-Oۃ�U�2�M��)�:���>�@΃*\6���+�r�i[��	>Ǥ��,��<����H1ԁ$**BJ�`�C����:o��ű059x�����M��*c�ø��ht�I�zSR�:+�(C�,�z`�äl����Lz{�}У�3������G��.S�"_��S�}ЖNnl-�xXý����]�3�3��+_�����4�M�a�n�[�Y���7~oDg@K�/�֐�l��Y�{0D#�0�n�7*�i�zn��%'P}!l�<E2#R��`���eu5�W1Y�%�u��� 5r��=('A	�dL�c����vf��7I�g���}����S��k�3�6����Pȯ����]���5�՛S��.�Q-��R��z+j1�RXlR�+a�����-��e���
^c�/��D�n�M���6A������{�L$V���@w�C!1z�ˆؠEZ��e��
�'j�}�PYA	m�)�uH�W�`Sb�{��[���{��:ld���6�|�DE�h���Vd؂4x��x8���(�~�\��3�m�o�_�n���.���������	�Q�1da�R��?Ү s��� �#��At��Z�	��100п�759��'�l`�t�c��q_̳z���QF��B��˩�_�Sp�j�3�+���p��Λ�^�9F���|��Y�	��o		�U짡��Jn�W�;����A��锤x�v�f�����Q�s���-��_�<+`Ǯ��&�Kׇ:�$��u{�޲+K�X�\��r�Ș#�rZ úg��<>�*RoQ͇�<?aY�p�;j5N�|��`�/ܓ��+g�K��LnNP�$��W�u��{#t��M�f��0��V���u���j1����66�&��>�$��7��>Q�$���L��.���WlʼMV����(B'�\MN�ϯ*)�BL�oqٙ%Xt!��^a��%Ի�{cz=�i'5�8�8��OS�L���S�꾹��_�?�xr��V���Q�v�	fh$W���<"��ԠJ�0[��!���%'��;Q�^g��I�3���ͮ5#z�Ւ'h�{�0�����F
�.�3����yHyV;�O�حsa�#���6��j����ig��y�[�����ZYb���{p�4������������V&fOx���Vև4��J9�d�LTj�W����8x�T?P5z�����W�A˖G<�������g�=�t�9?t���+�/����x�3�yE2�O#
|�6v@[ҀSd��{�8p��J�_���o[�a�F�u��;wS�K\����N���!,RV�:���B,H�=d>J�h���b�� �Eq=�tہ��\������h��q|xl/���93K�)���*���ͧ�.�.n�GKM�������1� ��O�!�
Ty*�1���γc���sS��RW�k�&�����r���<�2mR�K�o�/��E��ƽ����yG�����.���l�)n��T�� v�I�0�r����/��N'�q�0�
��[IS���4]苬�},��@�:�L.�ڃI/�O��R��zPqyI�/AJ�܇'cݺo��
�n��qP#Y�RBc�7���U7��_��� ��Ϯ^���m���4م>���(��y�gX�N�wÆ���:���!���)�c{B�xb;����e����,���̭�"*�H$���������FV��B�45��~�<��;��q�0��~��͍l�����K�౟���R�s^�d�=Z�B�O.<�Ι�q��:N�ʓ�k�nO�9$˛3(Rf,_��0�ݹ	��Ԥ����E����[/BQr>�Z�i�L'��|����{��x�6Pi|v�����z�s/p�~���V���������լ��(�5�>n����3���@r�ˈ�?#��F�W���a�f�깘�OZ\�W�bOoj�\GX�ט������|U���I��x5�4K�dt��	BuRl��h�lw"V�0�7�Z�Wt'lbM���s��!�t3D)��5uqyV�t����|�����~���p�x����ގ�O��������d� n���S `��ABW�����L�_H̃5����fK&�M�X�������]����7�\_�uTi?�$���yU��H�뉸~����N�u3+��-�i�X�Zn{Q6�[l�]�������ۼ��N��r���Ȯ��Ղت��uѹ�f���P����0=��3�8+6�}�z����󮕵u�z�o
|�>�"��C�`SA�>v_6�J0��J'����G�]ƶ�ͥ�^*��O�NE�v��2�h����٧�C7��^����ݞ�V���H���F٬�~6��Rf�^����9��6m!��nm�R*Ă�<�ϗi55�o[O����Ӊ?)$~�q7������sX9c۶��}-{rpCے)�4 d"��P�c�u���F�&�6�f���������s�v�ܬ^�В"HG�z�L�����7��g֩6��z��;Pln֘Ю��gW���+����d���r<��v��E��d1�,c�yӵE:���I��O���v�h�&��Dx��1��z�!��x6v�B���yO�Icf�&8݄*���X{���U�������@f��$�֔�С�)"*)�gK�b$��|��g�D�#;�'�����(A�,G�q�m�^Ǟ�R��t��suc�K�$��#������N�0w�<����e�0�g1�m^P)X��vZ+O���k|z	}�7�r�_SJjG�=\�F�C��{�W�V!��-Z�"Ts�Î�^��v�)���t��(������r��,�f)��;�\�H�`�Č��Y�	b���M'm���GiS��ب��B�>x$$/��� ͙�u�\���J��a2�f:|8�*T��W4OX��{�J�j\�?��U��|��ZƄ&����I"�_�Db�-��2�\������N�W�
��I�Ĺ�ܠ#�m��D�_Z��.f9�3�4�������>Az��g�&(ѿY�<!Q�)ܚ`�t�l}s���<�r
[����[][�e�765�h���I�	/:��w,%���R����^���)�!9o8��h1�@�_��}r���drke
�o��g�����S��)��{8c�S�B�h;}8�6^�38�]������i�/X� }e1��;\7@�r�#c:XE��~��lN��ŤN��ʷ�5}R���YFb0�4��+Z�`Mo�z2��ў��"�[FB�����pϾmJ���ͦ0���y�ݦ�&x�QMHW�#ڴ*����%���{�jwz�xa��8�2B�J9��iY<[�I�E��eo���׍0��)f�����G_[��p�����=�C�KY���fa�@n7�̓�[������5duZ��8��=�P.>>��tA&Fp@��hBR��͚��)��{b������.���r��s?Kď����j��KlΞDKX���n�,)n~��h�������f�~�4\7���p*M5aQy�̾���(�{8�w�\�_A#�����i����s�x�w��h��G�ɨ�n�9���k�-�Ѳ.��E�o@�Ǝy��_�~���.fT��;��3
c�d��^�Z��`&���8�j&'�8��?�b�w��Y����<g������pl��U�Q�|L�F��۪�<�FT�yJ�I���ә��9�i#�H|�����9_$���9Q�g��a4����è{�����	��Ui��O�P��������XIz�d�+�bV��h�b�t��?>�~*����^�e����(_��+�h8T�h"y��xK����4{Ȅ����ݞV��cO���K������fW��ݫ�
V�M������u�ڷZ���6�>t7yB\1G�6�^;z��d�Ơ����jό��k��?���>�}$�$�['a�������)�����|0^i�49�/[!�+�^��ϣ��*�_�������?(�����5(�[��5�c��ݘ���tǵڪ���>�W��ק���[�(u=�����$���+|�K�&�2��3��PL4�P�%��/�V�q]�VpP�
�.�N3�v���"�
}���AH>8j����9P!)vpN��,��ƿ
�?v�H^Y6y=z�Q�����"����lh�����ߍI������u��ް�n#�S:���Ʀ�ݿ�UNOMmx�����IӲ��8�	`͐M�[�rP5	�KG9��l��D��ʮ��倄����m�צ�Z�1���3GD����Z�4�g���dl�񈵃p"��ȣ�>]�K~��w799��v=^����f���e��B����M�SԷΡ�z<~�Y�ڇ�~:1����h[���4.�ƥ[^ة�׬f�����~�$�@�V5���S:0>K�+��o�W�UR	�X?\:ߩ�{q����tb{�D���C�T*Z�k]��5a��>��=I��oo>��� `�[T�F�j4�J&X�l2{��|�U�?A}'�g��Yo�|}r*~:7E��/�%����v�#ܝ�Od�N�h�_�����]|��s
صV�[����+���̶�*D����Uv�2�/�TQዿ����?� �����M�BF���kXsր����F�t��,fV���� �r�'6��=�Mq�4m�*�Ie����jܲ��v`��A����?KwY��}�C��H��Z�?��'p%~{w�u{m-��^�]�Od�|g;-�K�X]K%��o1OJh��'��D?KfD��i�|E��v͡Dua��=��%_~21oԾ��3������RF�Kxv?-Q/�&���f�r ��Mml]�cM,��f}�E�t	�ǋ�d9Q�����Ge셍)邾��fR�~�or��WU��PN>��^�Qc~�	���Rp�J����Ȃ��չ�w���m3�+1�����$��6W����G9�0��ps�*���-�O��Tڿř�*�;�ɳ��P�p�����:L��J�v����_���C���}yPh	��]�k*+*$�����\g:������4��p��>�R1w��M���(--�w2���%/ˇ�ձ�F勨�s����g;a9i�7�/W��~u�߯;b{L��g`��������f94�ż+[�,�cV���5A��1�⸕n������~��>�	Lh�,�VL�}��w�3���S�C��~�rO��r���pt�j��'<3Tӈ:��;}ۤ�A�,x(rf����?������h(ֈ�9�ݏk�v��o�5d���/	 ���ƖsK%��K��^M�B���+���[2��Y5倬����e�[�'a��"@��>�G��Lnmw��;Wr���tE�EvMZ��NK��N���@�8ua���
�%}^��r]*vݗ!i	
�ا^!<��K5eש�elݦ��S1^�gK�����<>�n��.����>Yӳq�����ַBb��j֤�TM!{ٲjZ�]H�v=��{q_�893D�[>o���+��p� �����pgraoq����+M#��|֥y�`�o�g�Ƥ�9?���.� ��~\L�O������������}쮑v��C�h�U�U]^!�����כ+��Һˋ��M�È9^V�e��P�ޥA)�4�S33boMס�ź��i?�?�=��7EP����K[�Q�o6`�Ӕ ~��L���U �4f��������)G�˯=.�y�7-�s��g��)i�}�;��S�Hp�DЛ�Ϳ!�k���N�u�q+C���Ķ�ģ�ºK /ڷ�߼;o�'�E�q�Q� /�y3�3=$[
Yp1�07��_�>s;2qw?���S��Qs����׽��3��02#��<������\	�q�)�b�G�>�W�>��<�}����)�D��b��"����?j���|�R�����[�MPp�I^�8��u:�е�bqH.vk��k�]{��^�:�j�a����CE�m "�����e��I�����$�9�}0��`eޗ9�v�)����e����+�	�2ڡ���!��Ѭ)/�k�a�c|uN�����mt_�8�����ɬf��5dŎ{mc�w]��5�S�^!'��x:��5���򶿷͸�֛�QV�Tꢕҭ�z��U�������pb�R�\n��J�2��S�jY�Br��M�-/b��mmq�yS�Z4�<�g�3�o���c����o>7�'����N���"��%L��������r0�N�߷)�'���PSD�,;��<�}��M�D�Q�� p��z!�\m���z,ђ��DE�Լ�T�qw��/A	A�O	�N����S�e����5��Q�fZC��C���� ��������̡�b���B^8����;6�<�O��}�߾��
�����*��֎K��q��\)o��4O[^���aM�I߈!4l�d��0���M��뒬��0�dn'
��:�~��<��Fo`ob�L�|n�m(�c���̇@ �y;On�]׎2c�T��lt/fu����y]b�K�c��oj�� d�d��h��՟�`[`%�~���=Qi��N�J���QWW��l�z�C�6�D{$� �s��V�?�m�j�<z(��N�)l����)%*+�I��X����գwY�7ь3v;gX�C;�i(�ձdy�,�X!�X�	I^6i:7K���?��� ۖ]����VL7�.��c�p����̚�2.j��v��5ޙ_��~ �����J�k���6c�ZnFd�G @6uD���6�XMU����L�ܸ��|�^��XR	�z�-����� R8x)��b��08�&h��oVQE�Ǫ�><��PV�?�@D ��xMe�O�s�%&`={'؉�A9��䯘F�Úa?;::>An�x���:|��M#�%8]�z����zR��������R�ƣ>���V/���?,��\��w���⒙�~{\��KJ�*	���c�;q\qt=~�O�A���m i@��ZS�@�\� t�`�����}����ppr�Z�<��O��z"�~�I�I௭J#��[���~����a����dP��-r�ЭiS�VSB]s��U#y����111-�灞�2�ЌT�"�w�%ͤY<�(uS�{�աd��= [S?Kn_1����|Vm�>��6o��×JF5_N������{|6��aɨ	�Y��5g��W������W'q{Q\���m��:������2[w�	<(�Xz��
��*F�'|�n�agF�6�[.g����Ҿ=Q� J�eV�?r��Q�-�xnȘllo���i��ٗ��S��no�q�-�LԾ��I��u�����1���t���y��//��{��~��?^�y
���G�jc��s*�o,�;�\�4��
"��T(Ѡ��Ɍ��DF�ĺ%�wY޽��/5Қ!�1.��Ǣ�2�����2�?�B�g�A/��2�Br[��|h]��"�k��^&W]��vbc�ι��"� �TnM�����&>��XE�
��Ȍ3���nP|�_Lk(�zSA9J����R�}�&�1k���B�*�OW�-9���<�]��{۫<)�%WJba��u�2��_�j�C9��*B�ʠ�����a�������1���nՒ���� ��$��?���b%ڂ7/L�Ű�J�~�jO2K���ɱ�&���z�Cu�K�Vo#��vc�0[�dM�<`�d�N�::�]?w[)�DM��{�*u]�fW| znYd��i՟�J2�*7��%Qн�%�JI�r�S��o�/M}�zk��n�׻���s�g؄��a�
�'g]x6$黸�|Wq�tt|��r7��ё�]M#�5c�ޢ�[�x��Zȯ���nZ��b��z�*�]�������%]��&�Et<{,$<�E�JR2v�S�<�ɔ"��i�L䓏:o`�m��%��*�&B{����D���0?V����{���mԒ-��dmp`���H1G)�$0�0�i��n���;'+eݴ��@�7�v���x)��gk��P�L
f������Ϗtn�&ud#x�Q	Q'�NL������!��C�O�-Ӓ���� U�������]K'S���2�8; �3���OAn�I��Ro�H@���+\���'��	oJ�{q��)�^Ǚd��R�v��3���k��̺Rp��w�=� mu:%��:z����1�T�k8x�X��bюʁ�~K���I#O���: ��0�\�'#��z��J�v���Y��C�;᜗��G���SG�� 
+x�q{���y����u�3�`�Dy�w���d�N�t�?����a~��t���$\�jfi�a\��pP9*�j�P=�,vp�޽�	5h`s�o��l5�9���{.���.,����m ��Do�+�]�%UZ5=�/*ި�iN�*D}�>*-.|��� #��T AY���d�	g{�l��J�A������M��Y�K0�b�W����A�۞-%J���ďA}hI����񣨁oB9"�J�u�4I;s�7��Lhg���i���� 4���?��/<פ.��g�ߪ.!�>ې��ub��1A|�W	h�I��b	���K���,Wo������If�s��j]a��m���7_E���!|(�t@�>���[$���T�(uf�t��}����{�>�%��+$��/�ڵB�8�4���?i�8GO��3�Ӓ1Z�q�E��4��4��3�_%���C������5Gj���l�D��wP8<9ꂇ�,�[��2�3i� c�`���mO�{:�A�啛�$���4h�Z�J�Wh2gqJ��(Z�OR�#���zX������j�w��U_q�!���=��t�N��S�?�,�i��w[jR���/'|���'Dfч��#�`�S�u{ǵ7��N���[ެ���N	���q����a�����NOS���p��\�q�*�J��Ѹ|GT@����$��z.�y���_��*=��s>�(��E��o�g�b�o}�ƕ�̱�3�H�榦���I�#��wv�e�%)�̻�J�8@��_]�(�7������ڋ�_'�����ѐ���t����F`A.#�`F>l��i���6*B!��K�v�K���;~�>�y>Q�cc\��ې��.��`x1��K�[-�~�ȣ�c�~>�G�+���)G�����R��R⽈GE�O�ɑ@B�����o#��̌<� )���-����kk�t��$}Dx����.h9(lTxO�9t�yxxF��Ի��?b����#�^���u؉�V ��c�%��1^i{�ǈ�L���A���r0[�jE:S��r&�,m���oi��ͫ/<�o;���r�������m�L��%��͉����d�@�Ƈ��j�!@:�E�>�]���L3¿���@E�4*ȇY_��`�iJz}J�A����2���c�^j�:=��W�+۪]5S�t[P�5z[�.�y_�'D�]�EW�E�!)�H2����_�"�j�d1�e�����[f��Wf�^��s�T/<V�3��'������s��n@��I�U�#�f�x�D�����{�S`$x���]�t�?���4����#�.�ݏ�X�_ňX���^ g�Z`M�m<,�����/Uf-��K����F��Se�}]Hֳ��XޒZvS��K�b2E۽ٖ��>I�B�4T|�O�_Y4�#�Fb��%v��>
j`n��_�ǀ�Ԇ^l��l�8裬����m,M��̈�87uJ��v/�=#/O�~5e?��QX<�nhږ���*R���ڤsg�]�;��9��A��~=��W�����%|��;`�9AA��Ę
!fڋ�p`l9�jTS���+}�#d��6�`���ЖL|�|���-��"��l���_L��Q�T��$��ˎ��TZ	�Q>Ŀ��x)�)�UTt�[��E�U�Mh�N;|�� V�s�4�&m���Y[��4u�.������h�U�	R5��97b%i���8���r�MIIy��vh~6����݆��HA��R�0I=����kc�VGQ˙���۔p+
<OOO��Kb	�~���
 |"���q��bp�����5~�	ЙK�z��V[AE����#�:�n�׌a�oc3�8����V�%��s��d�:���-
�}�ֆ��!��e&ژ��>�����3�sЧ�����8�-����(Y����ym��^u���fkt��Lf�?�XQ���k �~.�иƃ-�t��4"���\��6D-<^�Cs�Rs>M��h?�0�G�!V�Y��n�	�$�F9@�@p��6M �V+��?��~�o �*V�@�����g��J(ӴV�P����ػ
*�p~��]קގ��j����m^9Wֹ��{ƦJ^-ܖ��9���O�э��#� ~�l��KӦg6�{>=Qs�Ư���e)H��#O��p"�5�Tlђ�硴k�kj�#5Z��v^��8��6�MS�����7�!v�Gn��j�W]1m܆��&����d�&���"*��J�b���&8�i��A�t~�⦺�/_޷lj����o	R���Y���T��u<(�sy	��Y�Q�}�)X6�A�X�����,A%�AK�Ҋ�Htl���L�!�
iB��H�B��e�_�����Ҳ�9�ڽQ9��e��l����3�<TQ���8�&y̦��}W�" @H�ٓ�>NW�|u���x�K)�s	�����y᫏�� ?��E�W�<�pKħQE����Lo��?�g�Z��A~��S��'�%�W͢���ݚX��~ �(�M|"�1�N�i���,�����<����I��%-�|cJ[[�|B�<�^[1D���/߿_P� 	��m�'����W��e	�FG���P��^��>�,�:f��i^@�@�-�J����;��k���N�N�F�y����ϭת��Z�Q��MC�"�+G���ZC�ԇxa�.$ߓٙ����sߋ��1�������GK�yt�2x�X��;</@�icٷ��%�l�--���xo��1�Ƈ��jZIQ�?��9����7ʥ�&�\s@�@~x�~�^� �r��ʔz}���qW��K?F��=�)���+�X�K�Я7Yެ�x2�C�[ٟ>-/�Y����>�vm�L|~�v��~WcVSS+_m9���_���1_׍�$ʓ�]���OF'L�X�j�۳k��ު����T�������+ jCCx
�ʥ��X%⮽1f�0�@Ĕ\�[�܊����.�B���++�U��u���F�z��Z#?@�hT��;�8�>#e�)#�}�R�[�I_�si��/����K��Q~��]4�n�ǰ�n����ڷ�=b&tU�NM����&��-˱����fK�g�gj�T��Ѯ��2d�T���o#Tݨ�\���	��A�R�ٔ)�����/3�g��"$  �������.��z��RQs�Һ(Xb~�p���]wW-/��a>�ͨ����3���(�I�l�ǈΥ����3��z�f:??�˓�}��3��A����;4���L�p8-����D#����)������~KN����Eo����	�~�uW)�Z�1�kc����y :GFn���b����W�ڈ���f!��8�0��q�k� ����w]_o���X�Ue�z��ӧ���(���P$��t��,7bRŻ�]���6x��#�6�������p��kq/���U���62��!P!?F��~��vWu�[w��G������qq�j8�#\�ש���,%�����|m�*��o!�$
H%�n�e�ОhZC�`������f�J)�G��FQ��j��S8Sғ�W�3,8b;�A��n>��q��[!0�ae{0Cj~}$/�V���0��־���=�? L�&�)�.}5���bi�u� ��o:�����;YHV�
����h5���p&�:f�b�ϧT�,//󤕗Ӗx� ���dg�$s�	���c��ו,�
�,P�h��4T��Y1�)��L����������eI��j�dw��T/ώad�%��r�7q~N��{V
M�t���Gg��C�z|�Ͱ�n~mm�2��DK"����)�dP�-��!%�����.���xv��A�SA����'��p��2*GlW�Yw�����H�����Ϛڱ�庻�g�,�֌A?M��'��Ƣ ��)�纨(�3Ia_%A�q�|*�KM��&!h��t��k<�!�Ȫ��~����D��ϸT�y���:ؚ�٥��}�٣���*6�܇�t4$�!~�#�	�7o� �Z�t����z�����k�ð�/�>9Їz�i��"XK��8g�����hfb�������Erɜ�uݤv��u�3�@������k��@B�-MB����ʜ���%w�Q���/h:����yx�MT�X��|�|���R����<��[��sr���C�C�+�dXXlfd��ڎ'��[�|�*��X���7t6���yBrrrU��5�V��iq�l����.�`���y�PO��E��Bu���",&������>Sh�Fp���m+þ�=�o��.N6$nEx�	��q^;��� =���@�U��-M�P�����������J������3��t����6�JO$��ԡZ���͉RWg��&��>^h��d�Jff�wˬ q��]�9��s��5��m�Տ��Q.�;a��F{}��_������O���V�P!���n�����nX�d�F��^c5�|�dGT�N}D0�'��1h5<ߨb�>�w�aS���l���ɵ
�
5�Bp[�_@�I�.����������,ٓH��{k|���zbF�mkkk%��7x�S��Ȋ"<��C��sØ��v���s�<�ڜ�x��:�蚙�Ԑ�&�y�H���'�W �Q��h��C���8)R}�3;��u���D�)BY��a�'��h�-,�T�?��]A��~�$F9{��I�S��v�ZH��� d;�U(\-6�*�5�3����P�QX��&�IV��@�|���~���x��{#��ʯV�%Ȋ�����e��]�g��G$�;t�� ���s��cR��g����%T�;������JȦ���:��"�/�u5�iֹ=��c��h�g�3Y�	�}]S���}(-'g�okrO��/�>�)q��-� �!=�^D4�	��c6����n��� �>����!5\j��Sr��O�eP�v���6#o��R��7&zlpP�q�p�8m8
sHH͆`a���"�֖W����a��v�7@gi�-�k¢ȊuvK���5���Ʃ1�66�sXϷݍ�K���k9��^���K6���{ ^�Mq�6___��g����{.Pw����R���ђjL,,�U7
N~~-��a^��_�W�g�W�תq�w&)?�e��pv'���"=�y�j���@/��r_#��\���zA��jX�ܧ �
�J{4�ՔƗ"����:��?g;ڼ~t/�&�o�

J�-�)�<�sp(����*����R�#r�������}GTT��P�+�ט��@�7**��hC�y�^=,��xcw���-
�K8���vsK=�/ƹC��߈m{��_P�_�e1�|�˴WC�4Yu��43�7��Tn�)�}Ң<9ԘB��>�ߟ�@�h9�\^���\���l���t�N��@�7ǝr�h��s�� BR�CZ5�o�cL�)��;�F�l"��5����<�6G�Ź9]���voo��>x(9�E*�����.�Y��XS�56^>4��N�pf���^^�9"�c�\����.2����"���i��f��ˈ�|u����t).Y���	uO��1	���ɑI���C)��c9��1���ɘn���Xﱽ�Z��g�Jo|��Ch����O������:���׌����T�6$x�9�����l�"�j�G�cc���r�?;��tb^1�D�
��k�"M7��V)���>���.+��G��WB�S�5���� ��Z��	���]��j&��-[�F5�1�$��Yz,�������t�!&PbW����6Z3v9[�޲"pX]���]�>�mr�ňhA�C9u��k	�/4`�;���}�Rp��]0�q�*g	�,+Кz�6��<�ei���ӕ�M�I�rcjΈC����d=τ����Ǐ���M�S���r@8WV���vo ��aghh�T�45���E�G'��m7����n+b�$^�*��3$^�<�52r���p��\�"� V���j�1�]���bu���LzNM��{���v�,�I��^^Y������9�]�Br��u5��,r����n��&c�@`6ߎPǶD�:��h���I�a���N3���˳2�D� �B��gC��7-�k!R[5H���������-p�^��M'�4n�-�Q�ȒӢ@���u� ��&�j:���G]2�Ai��|DX��p���)��K�#��KL�Q�־�ug��q�����:�i�1-*�"���F^�q_8_� ��Q���~��t�=�?Ԙ���q>����ё����~p�@k�ޓk���,c��K�>����B�ƕ�:�rb_&�G��o����e1Io�<j�r��3�IȢ}Ǧv��_���_�޽D(� !����VS�4��j�)��j�g�*��a��K�7j7�OHη׶����㓒�TB���+mt:ކX^;��	�.X�=�D �u�zw��)��yh^ޫS�t��_@)^�>*"��p��b�����0AX�%�k���!��2,�5�y扖�ix EE����Ga�eY![�+�P�C����v�J$���&�O�cӀc���o�����'����}ٺ�`4��;�dڇ��v��x�F�� �x���a�L�k~�<-��O�4��J��7|0~��z�r5^jmP�|[ry�]�S�6,�~ߴ�\�9Z{E��|�2E��d(kzĽ��q���x�� }���t�N���^*H�W�DLB�^��e���p.I9D]�;f�E�=!Y���^./�{�܅��'^*jzz�ң��{PH� ��b�ŔA����N�d �������N-uH�u~�]�S�����:MG�i�N�{	"�T��%X8_�v�v+(����K~p���y��l�l�;��mr��p���Q�����̭�V����8����㇏����Ŏ�is�����m�YL7�K�y��¸^���FՃ+W��?z�?�7��<=�>8nW�$y�	�+ڜ��������}���)���ߞ�i��/kU�Z��yo,����iV�k�}��p���y/�N?t���悷��G�%�=�o�f�n����{��/.3#%��}�P`�+4�������y��dKv�������\sg�.}����w�z!����YW�<y����\���U�{��~ϧ�ǯ�KCh� +Z`fק��K��̎<�z�ҥW��7h C~랸z���2�Aj������g�7���s��-��;o������]�qήȣ&34.a�uK.�:M�y��������a�]���]���������w���Zs��!??Ƽyq�9�l�=�
s�5��m˛;�Y��q�̙����f������/o���goZ0#L ��<�����{��cv���]���9���e����L�<NR��d��`Q�9��u�e��m����2L�9�������Ƴu�j?���?{vu�Y;}P.sQh;�����w���W��ŋ�a��~~q��}~����d��h5Ao�� �]�������f��(��7m����^��5�O����'[����d��+���"���_�N��?��9�kkj�|�7o�������<�����i�S�4.M�e./%�%����tFU��m1�����?���#fOR8|y��
���8�0���[*�{0��o��5����~�ž;~����C��!vF@
����<٭�bRa⁗��O�8�ߢ�D�ךf"!�ǖ-_n�<�W�
�΀���}�z=��[	��E륤��nݿ���,a`cg��H���q�&mt�FKÂN>�J W�4=zԾO�m��,`�������xm�t��mѓ�����j��(xsc�6;�L�N[|��5�9f����ۖ�
)�����VvG� uȧ�	�(P�[�q��ՙ&R���������N�g!wz���B������p;����yo޾�����_���=����#P������ւ"�=y����{��N,*��Sbч�����|�V_�ni}%���G6��/y�Ƃ-������Q����>~���I9X$��b	��J�r�dVY�cyZ*��������������ރ��&�{V����߻>�4�j�������}]߿��{���p�~�8��.�r�.��߲���J�j=���s��^�����f����w�GYw�_�w�v��w�q���Th���L�+L��˥���J)��OO�k�$v)����'k�������gA{�Y	�)��w' e��$df��:��3��8�R5��d,2��&R�U�>!�n�l<zvރ
b��(?���j�lʴ1�.\�p�L�bM�h0ˋ]��cEρ�T�$2��΋��2��v"���Y��T6]q#�\��& ���l!���������+�͍�����/qJ�̛��.Mf����ѕ�����Z����L%�T1�sʀ9�g%���F'+�Q�yw�B!�X0OeN���'�,M��ߩ?��V��	߉_�A�1!���y��z�Cäig�����:`4��&�A�L���9��Y���3�����e�SB PK   ��X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   ��X�|�	  	  /   images/e1d4e862-170d-4bac-8b1a-e4319ef50e6b.png	���PNG

   IHDR   d   "   ��|%   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��h���O���&���1�T��]W6�GeJS
ҹtD���m�f���]�1��R�,�9FAA+���֊�2��DI)�6m�1�5���������\�{����������s��<��y�s��4�ڵ��X,�V�X�***����U�7ܗ���<===}�֭[���4�IN�:��;IH:333.�T��l��EȬ�W�7ܗ��Yk��ּ����_Zh��Ζ��.L�B��fw#&d�t��������ķ��������q]����^8::Z%O�r��/��Ύ�q�[!��l{Y���Oݽ{w������nrr҉��۷o�&b��P.�xo�	"#<55���R/�}D$<'w�f/���)���/w����ϋ�Ú�#"�$�|�r�E�{��D��i�ؗ PT=��g��Od�ח-[�B
��v��QWW�m�"����P�c bD�a��Aqq"�/_!Me���DU������92)�E �b���3c{�{M���������P@�I�ɧ��J�$�Ab8�%]џ����ا��ғb&�u`��[��=I��E�2��8���6����K�%��=)9)�O�(s�\���>3y�Br�����2dr�w%�}mOH�,i�8���6����ԥ���\�'#������v#����F����3A���Tz��;���w�� ΃�876;�ֆm��I#\�4AEZ���<#�Νs;v�0�ޕ����ܽ-�Smȥ�J)��댓LkF�|`|�{[������\��d�o�T�CaD��{��}�H5[&���l�g�u���C�n��k�p�Q[5 �H��Q�w6v5<<�A�3*޳r�JW[[�jjj����s�@w�`�8��N��  �W�Z�}'#�?���\��ې	�T� �!9m$m�,���\�~}�ڵ�7Ƴ����_�gƓ8Dp������,��񻾾�555y�GX�����իW��h�����h�s�6x�ӏq�TV�\�J��!Ni�>�㥀+��%���U/�Ѐ��xU�'oi�9�g���LoF9�}}}��͛nӦMn۶m��ٳnpp�ف��Q����x)��[��ׯ{Ě���]��l�3�ׯ����d�|Υ���2C����;/ٲI����N@�.9"�$g�ʋ�R�]F�\
�h�L��JXB/����������$���XhCCCNi�^���$�Hd�
��� ��9ق6R���2'��e��t�Nc�#B� [NI�@�E���O��P#�-Ƽ��,�e�w���$�����®?�;4��f�o=���b�A����	[�a>[��E�2~I��YW P��Y_X��I�a�n�rq���
^^u��8k�2�S���+W�T'�6\1�
SdX9�n�800���9� ����*^:���B��7%�K�%i�fF�b����AW"Fe��G��n���8��&�@��:�gN���%���IK.��8�l߾���	wX��o���I�����EI�ZEI�J���^�ڭ]��[L1]�׳7��u��Ϊ(�@�ӭ_�>���@�=��/h����)df$�.~��?��p�����k�yCA��@������7^�q=B02��#��Bi�B�a#d\�l�<�3��Ȕ�T��C�R@?�q�C��8x��L��aez�:;;�� �&7�� ��ԟws��u��ǣ�����?n,Bh�9h��Pz���*�;v�X�z�\��b�V���#D�3�Ȑ�>r?7!��u�t�hkD������	9z����ݻw��+"8�<��8#p�ԕ��4�`6���A6j�:�Y�~j�$�{E���]!(��}��yJɰ�sV�d#[�bD��#s���W��K�X��f5��� _��hߺu�wV
"�r�Ν;��w�?�x[��UL?�Lo�SO�e�h���/o�Mm�DyUu��>��[ѨwvR�p��?~���xe4�>t��ok'&�1�g��~�Ns��5SS�YoSM�W"�*x���C����EÞ=��{���������������������������n��K}6�xT����?�&'?z���3��ӧO�{����>�ש�=)+�\����W{{�'��{V����}_R�X�YB�X"�ȰDH�a��"�!E�%B������#�    IEND�B`�PK   �sX���F�� % /   images/e299bea7-de73-4651-8213-9be9a85bbb4e.pngT�X�]�: ����
�4H(�)���ҍ�4ҝ"-1 C7H�x��3�F.ƙ5k����D�(ɠ����@ t9Y�� �(߅� <�1��
��� ��)Q>����#d O�Hi��ٛ��9�����٭쬝M����,2�I@ *�����G�ޢ�ė���]yL$�xA�mV+�*��V�iv=�N5�P�F������Rlv���qE�[�NK&�����Lr�̯f�Az�)�ȯ��8��ÁM�-����h�
�à[?0Q��2���rٻ�1��顪y������}~� *����L>�C����.W��g"@��
+sJ�|.P��&ꕤY��yz�J";a"j��^4<�=�%E8^�J(U����>�?������23�+��_`�PBXX\�>�T����#���W��t�n�|��}�3�Y�������zu�hY���b�r+��>Î�뱱]\�H��
����we4��4��:���/����c��^H�~��)*Vu9��b��Zx���#�y|�F�ܒ
t7X���������uu5��zz���15���慓�p�[`2��wo�5uM�G�4,Kϵ�G�9��?������7G�h��бA��$��(�B4��Vf�`���9���GV��E/�7gԒC�N�1�Z�}��/���jHJ9�����ari�?P%(�����RB����T���7P3$ϼ�!�ʕ�6,E��Jw��t���0vsX�z��
���8xy�t�jgF�kU�_C��Jv�U}�X�Mx
�
D�7vh���(�N�M�x�����j�f�?��*��ޟ�!�7�I�6�i�-�mp���x�\�c�7^ɽ!��иR�71����/>�ʁ7\��l}�����K��`��M����7u��pY�[>{���RQs�X���?�4W������3.�>��F���� �Do���򶩔��z�5���P�R�f��ˆ��STM�!���%�;~w�So�C`wd�lb������kz�\
�5�1@�'��g��}(�0 ����s�z��Uw���R
}
П*��״t�U�
L��j�B��4_��k�R���7l}���56lx*z�������|��~s�G�\JTqJ8~4���yH+0�n��^�/0%E�#�W�̎K�Ɩ�l�'$����R�`��/~9Tp��Į��ˈ����߫���RR��[�q*�d����ܑ3��X��R՟�(���~��k��pG�r��I<��y�c'�5��K�@�����$��~KbO
�ur	��C-�'��|�-���'C��[�w5JgO���fk#9w�����s�R��Ϻ���^7��%�!��(����J�]�?	�bo/)oa��Z����f۟���SJLz��73	^�G��e�J|�1�p�l�r��d�r1����j�Awx���̉�����4X=��1��?�d��`���v��^W1������6~hK��L���a��>�axО��Rr���;��P���ǳ�����cx����>X]��z�������k'��;�nz�@�=�P��<���{6]���%���j/53�V�z0iWL��!�z�󎫫���
^az��-��O�)�s}袤z���ExWjLӌ\����Q4�Ϟ����q��v�!� Hƙ9�%��$�RDwm���Ǉ,))I��.6Ck�n\b���R"���͛��T�`�,O�����f�o߾=
|�]�]Ι��g�ގ�|ts����{t�	�V�${��wD��:�10^����[����?�gg�R���8��ʶ�(�M���􈈈~ZUS���wʈF����K{6��q�I�akI	Ryy���U�����vt,��c322�,,,&c+*؇����O��}wԎZ�(L@�9Y0u�k����w;�m|}g�O���ڷboll4��H��^�f�K���,l ���V>��'$d��<�Q�x�O���^���vT\/�6����r���G�c�����a�W;�5Զ!�9w�_A��А�J'L2Ic���5�Da��*,/��!��f���N����ER^�qm� �y(,~��u���^~~�ף���%�ӑ,VBu|򇍎�7�Y���Da�sFV��!��4xe|��,��
���d��p���$e��0���D��R._�p㳰I�Z0~WS���o��U{���b(����EUW�柦���l���F��lZu02l"�eo��b��>_��7�"96=�C��+�������İ��w?����Q42%��g����M� �s�(-���[j�3��t��v7~����8��K��[p�"���T�PW7�m�CqQ��v7�7��6>��8;}���Jq��o0�T�ŭ���5��G>%����4�y��U�"���a~/���ߺ��:�T��cL$]�-��Ѯ�X�<��M]G':�w�$lyQVFF��p�JTvzz���5��J��19"��
��M��}"RhV���3�J��Dn~Gq���`���v_J���d��1Cu;X�ҼM��G[f�d��_+�TF�%�3G�wFЛ�$H�x�~c�0�Y)���#,�7����/�¼E�}�����8����^g,)zd92,��;�g���L�%U{ݗcq$�,z���Z����zsj�i��4|�ï��h��j(�����%$����D�k��w}�Xt���h���55�{Km�g��#(n7"�a�5�]�)�Т�H�ܰ�'$ɵ��/:��\>-��\T�����YX&&&�dmDl�� L�T��c�5���:VB���v) Hқ�k��^<eQ��HS�l���R������hZ;o���[����3��喇@\�#5�#��;�Jz�ӗ��H��G���7��kn-ծ�ץ��O}5���&՝�8�����re¸g����V�Q<w��z�ś�ȂR�F1HZS���W-	�<TX��rbQ[zk#q�L�0��B$u-�R9�5���f���Z��7o��9�:�#��-�^�Ê�W�:j_Ą�o[��T����.���[��j�^"����m$�mq[��\7/���Gɜ�������x9�w���7� ^Ok�	�qr�j2�������Örr��i��+�G燾���N����I�ۧ6HS�ת_B]����Qغ��/���13c1H�Z(-��cX�Y�[VQ1ç��@�R�y�y�a?�a���@ߞ��+���U^�Bc�g]�Z���7�sXL �Aw�`�.鳵��,��؊Ʈ��v��χШ�Q��A� g�).�Zb�=H�\�I�57�8~�%��Tض�s_Go�<'mE����WG��NK�K[�t�H�u����
g�p�3�bb�FjO�!�J����Ȱ굞���h�'>��}���,\��%$��p���=XOt�M5[��O�
H��2��$ �EI�[H7�m�]#�AFʨ�	y��'�JV`p�e�_o�}2us�� ��zd�u9�VH:>4���ȀQʒ;=n�O.P�[�dz�����.�	����uK��t�tXZ}DT�'�܉x��$d�$����+�{V�p��ރ��:*�O��N�)&{a�̀���k��!��̱�WVt�o��7�	N��5<���ϰ"DS"���<;ZEC{��|8�A0&m4i҉�е����Fc�����I��:�|9/I��2��-����� <���]���}�[��0UT�bbc󋊤!�M_�2(_SR�1����� }*,���J)0BV�����%ءHw�O��v��\��@�P�&&T%]�Z����Zȏh�,D�}vf���'�+<���q6s����[[QEVPȕ���
��|?�\�9
��O��577:[*=E��<�X��Wg+KK�K���j.$���tB���gW;}�Xiǫ3=��w�2�����""�tυ�mg�����<��߃���f T-I9�o�d	:�_�59\�i��;�Df!��=�*>��2::��p�ݾ��O��^��W��A�>jjj�vĒ�7��޺�ʘ���s9O�@�m)F�9��
��U��+ʳb��S�����^0�	hX�B�* G�����"3\������\�onn& �b���ab��_�S�����{����沵�o���w���$�}�:Z9���9�2����� '2����+
 w%�	-�5�_��;NG?�6�eT»�4ũl=����ʾ��"uؤ����Z�(g_OGA���q�/kx�OX/����G��T�W�b[?�@y`f}�|I�E�ݍ�՞#����z?7>�X>���h6���=�(1����b�k���Yg�Xm�!4e۪qr�S��bp���]�3Q(3�m}�����vP��N���i�mfگ%��,��	�@���p����a���!���5E��ǿ�9��B'��I�D�{���㹮��wZ�3��V�t��S�a`����I��<��x�D7JR�mOSz�ˌ�`\D�~ ��E����j$�p{�x��m�C��V����� :y�A!z�r���Ϡ��χ�@q|[n���p	,BS�����N)юH�K�ǝ����c�����P�������,�G��t����՘�$�@��h������ڬ�Hdỳ���8!��g�#�����[�4:�x�#�Z�e��)Ό5���sD?i5�S�.��w�鲔$���Q}ot �fk-0%�ʤ˜N�ʑ�x�_��V2��x�O����5�� `�q_�\��{*��ڱ7љ���:v#s���A��H�a�7e�o'_o4�&V/�U5�23~S��4�DT1c�ww��A-F��z{����?xSH4�`!� !D4�U����S��{VO�A���4l�����o�WNp �`�( ��IY�0��(��c�����&ڂ��+�����)i%�������w�|_�A�=q^�9���k�V�Q7,���?�1�g������R��� g�vE)V��鸚��@��q5��t� mط�V�@Ĳ���v�����h�v����@`Ƀ�y.�"BB�@ԭw���H5f���m<�1�<w�rI������3G� 5Lbt<Xxe :�z���Iz7^��&�-��ab�BU=���t�J'�zv��<+K�5�����[�� x]a�+�^<q������vh���͘�_2�of����䞫O։�R׿�G�����q@Dc>2[[6mmm5�$�j�Xi.�I b�./%4��U�9����w>z(. �����U�]|n�7�� t�6 ���|%5~�Ex�V�w:P-�W9o�D����H��O�yv�$�P�@P͟��x��H����0���;��!"ȣM?�˗|��<�C>ä.q�vt����W����Y����fk$Zx �F�.�������vՁH�ڔ�!l�y��2*�_K�[5��$�~sٺ����j�͍� 4����1��B/J��Q�p"=�z+GB5.c�?�J�Y��lۧX�H��������:�u0��6���&N��Kܡ���5)v[ &j[D�a�GX�Wk��
jctLg�����|�(�$��?�����56�hi�O�����U���pL���A��-�HEZE���&Z�� Y,�>�>*c˯��V�^��y2��;����$��J��1E�Z��͵��;�.�1��VpW=�p��f���)a���OB���%�Bs�|��(��"��a0���G�{�����=	lpz ;#֯�,��������?�c]��16#z�yp�8[�\?v�w����߃�"�Z�}�^� )����J��?�#�OH�)�hG��4A�ga�EVD$$�@��F	=�� JܚZ�fs2.(�8�C�*�~�d�3��ǈcA~�Co�ѻ�VW7���uL?�%�6�#ݛJ'tgGH�;���AYwwi�����%>w�t��g�Go���2R�G��
�u%P]@���lnF���m|�&z�ɸz�e(C/�ӟ~�Պ�NN��9��4.��|s^I-E�x{Ӂ�6�Cj��o�����j:�sY6���:�J�^E	{��=�pޡ�����}�X��g�z�S+��Q��׌=Q�T2@g��&���la��(����	g��ζ���30�ɯ��f��
S?K!&%�YOj����c�8\\&冘��>z��tB��wk�ֽ���:sI��Fk�Ds�"��d� ��~�����"�f���G�H�%������hLј�0�+���	U�3���04J�K�����1<W��5�x*m�S� �vr�H~p��Yj?O?��`݄~=@�A�iy]\��U�����y�A1<)��c�N�l&۔җ6w��.�0i)�9��.��$(�1'�(zô�U�H��ڡG�#R>�
��rO딲���&z�2���y\l���c$|-�l�9h��n[y����]j�BP��sP	�o��h>�f&�_�T�n��lW��"��V\�Ԧ�'÷o����X���)�e6fk6�C���@�8�pbA��i6,�Y��������&G9�yն#AE�k��G�<�t�SZ�Pɗo��;ȃ/����$&(3�_��
������>�y����㚁b��x[�l�;�S�L0vuj�s"'��x�"!�Q1�|��#j��m'ڒ+��r����
^2�HT��I}u�O��PK��-��Yǃ@��D��J
{�#^	ɲ��n�>��:�_l
}�~9^�٘K�����6���x8V�>XQ� M�:��l�G�RZ�?�u������}�\>�iM�Qb�\_��T lƤ11��l�-_A9c镄�����)+㪶��<�Z����Fkrb���ab�w�3}����;(%�M����v)&RěszF1щ�=�
P�`o�A���+�pG�!�Y�\x��єZ��������}���4����]O@����xz���PT��c4Yc�ȵ�bU�k�D�[[�#�$o!��83RR���hg��������|�y�%����n�c"���b�=�`0V�w��#��6}K�y�p����(�D6&&���{���'l�����EB�e]=,ZD��ص�Y�3����K}/��%�ю@���(��r��58�Q(�,�Xl/�~���i��0����RR���
�D׷��,�W-Ӽ����9*^~�"A0^��)ϟ)O�!!�ݝ��팁���	�����]'�&�_�������c4G��U#%_�|$;��+IӀLb�H�^w
�_C�������kq�9��]�
��K612��V0uh��7>Wh�1�����0�v�";��v�I~Ƽ>h�A�����4(@1�?���fבOQ�J�ob��GJԹ���,��#��3抉�7qs#����a�Yu�km%�PƷ����Qklj
�ZZZ��t���j�^>�|  ~��j~��~iii�C��ۿ�]\]���@ :�nt�6:����'��|G>�]Lc�j '��% �HHH ��i�p��v�^P��=W�<:��2G��
U{�����;/�X�h
̪�����euZf���%f�.rh�	nӢ72b��(�U��q�l�.IX?k�
�[�%�_h|弉֪�Qo;VTĐ�0�U	fnniq�>��v�ӭS|�lDP!Ui�l3$Y��FW�jCccb��z��!���lğ?���ɝ� ��� �b��..FH���]H��ܟ=+��A����j��]KEGghc��ӱYvv6too؝Y��u���9��v)(/G/,,D
������] :��t�JŸ���WBw��]�yNO�HIe%b�3 ���ք��i#G%�U�_4�=�&�;�������Q"�/l��ɔ;�/"�B�YZ���ǽY�>o@o�ǜ��`q��6��f3��z�O�����S�&(��ڵ_�HvC��w lV/��e\������,"I�ܜ\���c�P9������)`/��|��"*q9Є���#�\�b�6��}7i
��F�������Y�*��q�qx�tY�+8"�� ��Gԛ�D�j.�s����i�A!V�}$�N2�u)������ c���FR��@�w�! ��^
�xd'��C�D�zV��@Ai4�zkX���el�������rr|��JJ��?�� Ve��༞�Qn*�>�D�-#���Uf1ǪZv%I�������"�	�E"�m�A?��հ;óV&(�]M!��x{-ubR\ML���1�Ym�\&"���z*���B+�
��o�O��_x�5g��]��>���N�r���W[�x��D��i~V/�O^�]�s�O���2�?c%�m�U�`���є%f�����r�4���MwxLO�ip�	k�d��>�Ig���u���|^ׂ��!Z��\��+#��J���u�����pt��*."�N,~sNրE��x�����-I$�"�_����k���U����|��.��ٿ�3^�H
n�_��9O]ER5h�٣��i�/5i��Q������t3���I��{�ؠ������~4�٫7ִ�Ɋ%<ғNɤ%��o��A�5ť�쾥T�`�@.�./@pb!TXR�rat���߱����b��g�7萰��:�E��B�2��z�ə	����īZT�QG����V;�0gnS#�ur��'���qѕ/���������}�.���D�RŖgR�d���8�"[|�E�R�!�iS'U������łG6���M�h:c��<����(j�r>\�L��x�����6�{JR�x��	L �!AAڙ?{�%�O�<"�KSZl��kq�eP?�ٟ��!�W�\d�S�Vȴ��o/5��k�XÔ��9a�2a��:}���Z�����x���ɪ�l�U�����Y8555�����H�b�N^�$G�Dl:\U�Od�����k��:�e9�%`)�Ĩ���RKx�:�A��S!�Ѩ�x��?֠Z��/���9��.х���s�0k�`?�����	�6�&��R�a
y��;�H'���SKm!����y��ܫa���tr8����UW;�[�olt&І�m淒�����`�F�w,�����0G׉�M�!.������}�Rh(�WP:;m��ҡ���$^�V�K	��|�MԛT���c�2%\�z�%�+�����z$��=�������+��h�UZ��F���R�MGG�i�M@�\%���%~G[����$Ac:�	/�
�mE|2OK�B��h����R��H�x/�/2,�w~5𕉹;�ª�l��
���.�2T��4'
<�a�ƾ���
�Q���sca�ЪJvS��}������71�;��(�wƷ�Xq
�9H]��CzG�n�p>��0	�߳K�L��V�쨗*��:�ޡ���n@���,�XF��LN�s�\�?�%�uu�n��J�vOO���	�X��]��vd7t>�38�A0�`i(B����ې��ߐ��.Vd�9E���B �=Ү��LҚ}��c��c-��C
��Ib���ԾΪ�� ���@��y#ʮ�G�5��&�A�R?��;$�`rt�����*��N�)eS��T{`�M��6�T��a��pP����v�קo�0�6b"G6�K��}�>	�-�|��
���ę𺡳D��`0XE�Cʌ�.n��(�Ȫ��LLOo?B�صH�ꠥȢdz#���u@Es�Z��`����3h��e�0q^�$���k�_C;Rb/~!�����O�u���B�����F�A2^E)NA��B�27_���0��H�q��
"έx�r���oULj�����#/���X��l�f�~q�OF��4�4Ͱ�"�$�!m�TYP��V���Ms^�{�wN�p�:��䌤����u��b��}���ed&�z|
cC񤺾��)(�uW畗ó�:�͂�GX��'^�3-#]ǋ��m��(�5蟺��� `�x �e�͖|L��`-�� �%��KM=DO�^\�b�	��B�ԏCa�7=�o,ŷj��6K��"O��,ᐹqɌ�a>��B���A��>%�
13)�,D�	����h	P�~o��*J�2Ԋ�F����%8U���DI�p��� ֎�R)UI*�ޟP"f�_�Y���C�d�4�	��C����7�m�a����<k9��Nn�b͹�W\����X"���w>Y�jh������`I>�o���Kigy\��$��VǊR嶀�%�F���E�SgA�08�?(�Cq�r8d��z��.Z�`�Ą*&f��e��z?i=5N�ʿ��|O�Nuw8.׸՟� ~7t��=�"j�q���w|a�n���Y6�%��fC���yԭ
zj�kbV���/�U� l��[�!*�Te�u/�ـ�&]�$LWIF�֞�<am-�`�#� ˥q���C�7 �K_*(+Rď�.�����\u�Di��iF��A��P\̜pL�>mN�� R��of��W������������aА���������01İ�l,m�j��,�|��{��"X�c�˒	V�z�229�9ޝƷ,�=�=��	��(n����+��=��h^��\||�e�Qwޗ�H���'F��x����T�:=���HT�A;W7�^_�z��׎��*�Lje1r%��13�̫�i��o�Τ�P!�~��,:���jxf~|V��@���U��)Ϫ<����~�r��Vr:�e�I��L��Z�֨o�K�|���l�-*B'/o������0�Y��;:���*�7��trA@1�`%��#k?@=?C9۶R�'�w[�d��pph8߄��3>z�˘nQ�B+e�yTC�oo��� )T`��KO�
) ��ubv�5��(�����V���L��Y�����"�j��F���+��8������ru�A-
m��k�fPPRZ�EE
�))/���k��N˴.-y���"��ɭഩ��48��%UmvfL.S"�H�꽒75;�:�e<S�<�$����e��7(d��i��j��� �e^���a�y��{S0E���$��b���0�v��������FCp�i���iA�AN��T�,��R-�vY�N
O��w�K��G�f//Um���ײ��J�a�	�@ZU�;۝ց̢%à��5�u�����^�E���q��}X$�t��^]������@'�д(�GK��P������uY�$��^��f��F�
��U�G���`�_��ML��$&_�x@̢O��j]��V[\��ZԤ~�b�;S.Ϯ'ǀ�� K��� H��
������B��������8�͆\�q~�-�(��"	�CM��z ;����#q����I�l��@8Α()e�
{��2�F���������$M���q�L�����fJ���cLLL^G%P��XF�8�;�ɤ$�`˻E&<M�֟ ���v�(�	^~�	is�W��VF&���ʥ�����|tzz��)l�Jm{U�l�^���d�{c��B���m:$?��z����N��T+�>�Yq���֓L�˥}׃9RX���U��^m�#T �@�	b�k��O�-�Q)o�����5��+nj�-����H�xޏ����CK�1}�G7>�Y�����oӵ�s�f�z�mpX���{�٥�P}��""�H�E�_�}�,�I��V�B�dw0R�!n����4�y-���bIi�`��4>��I�u
ejni���V�ӈ����z3*Z�Պp�~9\]�].�`[!;F��R�F*-���TI�5j �����]���T��|�X��m�(�~ܐ]��fݏ�5���9c�݈<ë˽�;��H�M��ɔ,~���
F�4vp�����-]���-�g5�ɡI���:�,}����I�VT��y��H�0�V��P
Ђ~9�t�ii=;�Q��"���@�c�gf� l��1Ž)M��p����j9�is����.l)xП��b?=�+��TLGGGzd��:�\V�����Cqv~.�b��܀h1�-s��d��4�eK��RYȜ���!�����q�jR��Dd$������5� $E($ĵ~ڵ�VXP K1�;6o��K�u�ԫ~V��Mj��6��*�#��,�F&�x���0W9%|��_���
Op��R�F���8h�Z��\��R��A�	\3��3��Z�NR�޹d�F��=p<�ܴm�_�;99!�h�TU�vۛ4xf�c����СH3VV��F��Ӭ9}:��H$����L����u�����Iޟ51�C��m��	K�BZZ��H2���zd[[[&���Îx����-[8���lޠqI���D�2�D��:�&�Bg���a���RW�oo�Y����ƀ��Gڃ��r=�����d��9�@=Ք���%�V-m�ת�_*�ʋ�\����W�r���_�-F9��^�[}	680�����Y�`��FI�9K�h�����Y�������~w���x�,�U����	U<j9��v����[e���c��j��a�)��/�<�0�t샊� 2:��}Y��
d	�2�I��45�ү$lq?��8_�k �.؊�};�^b��s��UI��0ttK{�P:9g\�n]c�����]�D_{��!T"cu�1�wvV󗵍��0|��+�����K2b�����lv8/^ݯN�ڒ�v��/��q���'h�	�p�����$L��{��u�C�	+u�Ī�%��~��33�0�!9�;۔�_c�t����d�<��T]�����z�L��������L���VkV9o)����|�d���z2���ρ0�^=I�]��D5�R� *<#ccبĹ����V§�<�����J�<�S�bڹ�58�2���Be����p'���i��w���C��7PE�
��=��?�򝯗���đ����o��d+m�g4�F˺ſ8�:�p�oki4�ko����!����F��?�����TD��OD`b�X�p�?}ç��QҤ4��%�%S�D��@@����Sě�@�x�
��}(2<<lh�Ͳ�ʋWDFu��`���,.)�E���J���n�VO�z�=0W�VC���N���M� * 호�]������:�ۙ5�\�(h�7C���T4$�)�}�f/�,�>����HjT�D�#��z��<ޛ*��/9ЦE
�S�5��Y~��:P�L{vh�r��zlZN�4wz��H��#��@�4ް�P���xB�0毡!U}���D�F]��Ń+�/����t8M�6TXo��:���ns,�J�Bhy^�o�N�[[�4�� �9�Ɗ��F+?�!���:�E�I@�kߖn=��qH���d�qi�y/߼��{�7��f��?�LP�?a�2gv�h6b��X�:���ɺ\�w���t��Ճ��X��Cܗ}	wP���p��-��F�rN���/r\ �HAI	d�l�ӏ��&bB}��,x�j�E|�����Vi�MdGDX��⏉T��I���^,Fonn^ݵhŗ�����:;A��0�w��/���<h��>9AE ��f��<5�dF���r�4_o'v8�k�N�j��Ic��Q�YO��1���"HT��yC�M!�7�����]�g�8� ��qr Ϸ���_�̜κ���B��$p����%�Y�{����W�������"�`mf'�|���ͨn�'����"������
�肈����i#m��C�?�ﲦ���/W���DJ�roDj***�H�9�:5�/,Č�*y�QX��rz^��#ugm�1J�2�G���Ƅ��{�q�tx��W�_�=E��O�E�YnN��o�e%�[Ee��f�ů�eo��bWxr��/�VV�k�j�R�f�6 ��u���}�w��3��Ĳ���h�F?ث�:@r�!aa.nn��ѳsԐE4VAm��qU�ϒ&�eO#��"0�Z��N%z�� �<h�����ՠ٧���		�p�b6������aqR�AZ8�Uf�X������Q�Ӡ�8�I��e�����Y��L�piٞ�A0���Dg9hM~��襵�����I�,Q�7�sô��a_K�˟.�YW�aiJ|��i�0M�:՛�ܓfS������r@�zW�mr��
�V�/[���d��9P������!����	�W?�MFR*Ci!Q{c*@{|��G��z�5�!>&���}y��H΋#���0i�� �(K����նn��u3ID``2�>Ѻ����d��@��Q�\4z_��&�Q
3�Z�}���"1�(���x=;\M�"�/5�Œ�ٲ��)*����ݎ:�N`��]��&D]�-!�[$vv�6"G�-ܛNLs��א�U�!����ß���ʶ���|�BMO�.��`��xbآt�X�;j(��w�ʇa�ǎ�6���F�c�T��)>!໒O8r��PGE��V8Hm))���ill����߅îZ5�i�K]�$1<��A����B���mۅ�VJ�ς�A��1��b����?��W7�\>���5cZ�v���]��mX)�C��G"����t�j�3�� Ґ��A�X~�v)��0�}E/���GDL��)��LJL�-K`1FHHXX��wHP�FOP��2�<��e��	�Y�d��)\���ڵ�����x����^�u�XP;#���Jd���eµ���=.��Q��h����& �_u��i�Ơ�t���-?���_� �3ёuiR��Ƒ���I�t{��Eߌ�(�lERTT�FγL�З+1+��ng�H�t�!�������n�O�J�
��xqag�� Q��T�w��te@T���"\u��crjJJ� ��G;ֳ��º:�찲�y�n"M>W'|�ͦ�#Ӆ,dC%�+TE�7����#��:�|�]���<&J�T��s�L���(py��b��9=��l��ժ��A�A+m$�!��	D\���P����>� 1(g��nT�[��L��Ċ��?�ɉ�W ��59�m���֫J$��5���SP�Q�O2}:[rY�c0yI��/�p^��N���!�utL�M9w�>��������zx4ݴlb)� G]��s�<L��ڪ��N�þkwi��V������k��ݡ�ct`÷��	ǟN�P�
����/��,��NEùyj�ͽ���b����U6�Qr��f�0�n�E����yޱ㢢��/�at&� ���8������� 0�ˋ��ߘ�5��j�]�1оq7D9Q�a�L���9][3VPT26�,�A�MY+
��J�ɣY1�,��3m��$�c���s�;��MK�r������Y/���Bd"�?��M��ϕ��1*��`����)��u�)�� ��z�	��	�P�F��6��e���#0w:��M[4�*RWO�O�$��üU�޺̭��F��DO�SQ�����a��t�aC�T)�E��.�����a#3���S�j"e�EF�J�c�.x7B�qEy��}�­�L,�-�F�;�:�V�C�x�k%��_;B�ll*�~1��u3��]P������>��ZEFF�9�F�W>Z`�ޭ��������LQ����A�&�$���֨J����^]��y���y-zJ�A��P��"�U��P��N�n�^��=G�H]�b�~a$N��Ǔ,����+ʌ��� q�t��ܖ�q0�������j^!���]�x���k[*�c
ǟ�2��휖�dq@���;�s����d6��W��9`��	��Z_!��v���˂��W�~,�9N)uy��~�@�����jx�zA�D�&�e��y�F���w
8t<ɘq�*3]	����`��S���$���k�������X��0˽{��$ņ,�aM�c6���v��=}B���9�&�O��5{�eOƨ�������({_��QmZ_}T�}�'J	��ML:?��_%���$ph��/�X 0����އ� qU�V�V�#��l�ɝa{E�����/5:&�/z�'���,FS��V����ӾΉ��jV��>f��GB��ޮ��D���˿�׉����w�Ac��;2���-5(�sȈa@�u�ʩP���4���-P^)dI��uvX���:۹o���R6���G���%���_.�[�[��\��ŹYE;�C�Q�Mmb,�Rf=�fשl�3�,��lLHLM��:�dRf~gz�++[/;����ж���H�Ӻ���{� ���1�`��u?zHf_��o�S�˗���â�.���K4�%-=��C���|�v�EЫ��X���IF�g;���Hs����������[�6��G����_V:�d<�xP�|O<��$#Z����#�������gk�V������JH4dwqrz�|&��^��ι.�Ҽc^�k�~�Z���+���oʦQ�C��#~�ϯA��s��z�{C�G8�?kT�S��'�S1<��^���,)�	3e������W�}�k0����S�t�AT�,�V��b�������m[�;�P�/�
\�G��7U-�����m�x�2���Ӯ*��B�_��v�2�|Y�gZ�o��Ĉ)��ܒ�fn���eN�w��N篔C�0�LM��g+�)���m��NP
;n�z;n�hܿ��p3��5������l�9�0�.�4q��h�����dr/)ͳ7���<
Ea�bEՃ����=�}�������X�}�=6V�r�|�=���M�=�j3��I:h4���]d7ѓ�k�`m�dU_��a�¢"se�ˬ1�X�D��1��*��o:i��n����t"����nBΌL��ߩU�Ҳ~�ަ���n}���,ǔ�J+#��%��1��8��R�֚��m9��&��zY*[k�L�^����W��@L��,��I��D~-$����X�)г����֫��� ���b﹊IW(��zT}�E}��`�[N��m���C�w���EmI$j=j�D�5� ��(Ct��A�&D�=F��f��Mt����{�����������\s���^k�����L��'f�>b�Rq�]^�4su�+��#�===T�������L��ȴ�q���M1[�@|�ΤJ���eg~#�!�ٹ��rq���Y��].�s��óܦAO�]���
�l����	�AL�/�
9g\�UZ�?|��ͭ�J������`f�B����CDD��Bzp��6����R(��p�wE����!�O�&�!��	�΀a�����rS��4'���/��'twL3(�U,w��0~g�;�7�Z���س���r��Ӳe�z�R]uO��9}|q�����D��<9���O	V^���Ku��C�:��(H$;T�`5���l��r���:�8z��:44&������څ@<��� ����s^��J{���G��2;֌��C�wll̘�BE��32. �e~�@ ��;0�疔��ޖ;>k����L�WF��+�!]�	��=J�����LZ��ϵ��֯QU��0���K�`pj�j��LF:����Y��Mx
��#=�7�d}v��5_�e�Uj~Ƽ��C��~�� 	�-$-��343w8kG��c�=�Έ���dދ"u�1�t0�͔��D�w�R�꿲w�(�g�>fbZʓ���-��|LG����ꩶ�x�����}z��g-�_��a��]�^��B�t�]j�Q��S��,�mj�ħܵ%%݇G�0(�U��K^�p������q$�N��'`?�yyVq� �[��h�E-���6����yQKb:/��;���zIڤ�3Hh>gj1Di'���a<<32��yeyo�ws�������|�d������K��:�>z��T�}��!t�Ь8�W����́Ajg6/��s-����A����$[����X���tiX���#,<5�/If�6��Ȅi��S���4����v�!�O2��a>ą#������3{!���d��~��7lmmY3d$��l�mUb*�3�����9�Dի9&7,�[�B>�m�>:y��^X4#���!t���4�	�J��0�(��rS����/:�І7hh'vw1O�s�4z%'�X�Q�Fv��,��g!q9&��S��{o�O�Ʃ�R�W�
˛����P3����'��0}5%)=ÿv�W���r  ޺+'(%�{p LI�{����ʍ���Imq�UUfnj��r��ç*9jGC���H�_l"�0ڊ�E-q����+x�����A ̓�[jW|��$�.��'��'��A����J�����M9�}Y����ͧ/�f�k�>����J�ii-\\~-�z'z�����Jib�r��߽��)i��r���H�R����z�3 �����}$L�㧍/�jP.�$�5�p�7�]v}�
G�y��6��~ǭ�1�1�z|�߂�N|�P�؝���L��QH�%�Pe+Jq��ͅ@wތ�?�+�'�������;��K��$��J]A�Hl��O�Ӡ����E����?{Y�C'�������*LB�M�ޡE�S��=`6��5�c���z��X^�xrs���pĨ����I\�+˩j>�$T�HqA)fm��6�q���b�¿&��$<�=)���7�:�������TR�J���� ^����A�9�x>��g��|�}IOU��7;��C��նw��+2���C+�4�|���:�;k�X|{(sƉ��l�J������{9��wdFQ��6�[j��;��´E�1��}}<a��. b���9�xt�6ة�k�5�J��^�D�	^ɭ� ��������?0�>���Y�3�t��[�3IIO��j�[�-扚�P���^g�V3��r��z�7�O���^�x���6�v�I�4���bH$AvW�x������,�Y�]�ޯ&���{~�H�~�����g��荍*KEw���C��r;w�cP�:r̖�W�I��vѝ�<�x�y�`��@9���'}�ڣn�h�%���|�&���}��P�5"���v�q�Ds�u�r��d�LR��Y�F*����}T&H�) ���:�u�6"e���~s@U�JIm��X��C�v�"�G����-+�kEs����	�+l��@���KuJ~mfQO����]�;pL/����CL��6맽����{�J��f=^&�	�b�_L���4�jWϒ�O�F|Oo���~����c�<BL<`��?�h#�a�q��drP�E�J<$��bQ���z��NBW9��j�k&�h׸��pٝW0�[+
?�'�����_���~-O6�{~�j��.�����lʝ��6t�������%?g�t�*�|��������4���\�w���J��p���$�)'͍$���D�q��Rpk�+����<��`�0��$��2#.���V;DJ <�\����W�
�{>�G�/gfؐo�lnnNy�{�2�!����ʍ���g 8>���ه��y��Ai��oJd�~��B�E|�|�2������C�ח߯��4��5�\��t4��W��!����� `il�����G��)��r���ק[���0�b�=�=c8Hl�[ɬ����R����\9e�	���gd�$�$V�ȝ�ݏ���V����l��"�a����®& �UWt���ʐ���dv����g���A�q�R����H[+�S�Կ��� �C`&�?��֭5gWZ�f�-�fƦ�3���*�+C�TRh��Z?�o�� �v��`�>��mEC�o�y�C�v�](�g?m�� j� ��S�XB#{Pc����j���r�w�44��aŧM�	�Ǌ�X���'�ɝ����(�
��r��@���d�a���/q  OO��(Սjm}��~*�熛�y��o%�{p�+i��I��Nk^kF�k���Pƫ'���PRO--���Q
�Ư��斖�O,�?����#c|��ne� �iӛ�3�OV��esk>�~���$�o~�Ծ�Q�]I��.7$ �
��?<c��G�����[���Q���z�l�����
ź�j�ڤ&�E��:��}����/G:�g��� ��q� #y<�χ5�}]AH9��N�|����%���%�ͯj���	�~.�ǒ��Q��i��b\�=	�	��g%{v�fdl�{x�Hi�3����]'���=� ��^ɐ�n��G�������ѵ"��:yx�!���E:;�m]\�������.����������?^��B�L2R۽OJ4;M�����y��.˓����&

ZC��n��/ ���_~��^��>,#x��5�(ڋ�v������x%�S���%�<!@�ug��;�l����a����=��] U��û�X����i�LmD��$�.Ŀ�D��'�V]ܧ9�5CUU:�-�N��b��J�SE��
���fN��_�����\��G���?UΨ?6n�*�@�#� �̋�a�WJ�K���Y�8F�W5?c^��bǻ������
�f�4Ո�a-0�Qq>�滕`�C�z�����
���Gtg��N���D-]:���Y����� ��}v��0 RWR͸7Ȣ���i���p���wZC^g��UWX0��@�[SmG�߾i�����3u�q6��6FS|�y[��ޛ���X�(�Ҹ7�%!��)RLT/鶩��E,0S�����������U*�lbX���4�g�����̶��Ϲ�k����o��4?[@�S@��9JԽ���2�� O�஝��xv^�t�h@��1�?C��9����B6�0�E$�֔>ERjFѺ���,0}#\�~M�5'K��
�����uh�?�B�39�"�<�d���������,/54H!&N�t�Y��g�ѩQ�H��� �~��s����H�$��[�h����v�3xr�IL�{'�(k�L��9s�Ւ˗����C��q/�댦�>�l�B���dId��=4�h���4Qٓ���f�rq�55|kb�y���8�+bg�!�x��!+�-�%Z	�d�[��K�o��P1���\��	X��8u�����l�/BZԶ�y(�����$?��l�1>2�eB�xi�7g�zV�<	���CP�,�`�d�����P��[���tP�Fw��KJJ���_����Y&''�f��r�oFǃ1�Gk�yͶ�=����Y7H�}ů>���r[J�a�d`��kk���y���S�I�N�	�\ρ��mll|v;�K�,�����1O�rww'""��ہI$��ǲ�R���F��Е)Ws^�G��(Q�RU]}���/l�=|���>_URx���Wh�����0Fo�z�5����<V�0��EP��ͅ�S�X`%(m������\���c��� ����lN��e�����d�,�����_��f_Urtb�C|��"&��%+��zO�A�Ͻ�Z�H���h���	h��/�@����zI�k����~����I��.q��酶Iw՗���`���?>�{vX����Q�@񞛴��P�H>sj.� �23��ڥ���v����XF�h���e 
�2@�r[�
�;/���RB�Wĳ� ��J�gʞѯ������z����oo1�|!�'�Ȝ���#i�%�8��-Z�y������&�@2t��\N:��u����M߮�}�����gs.����M�S��'w��ӣ��Ўś��b�=����L.�Ѧ�����9���T�.��R����$@�UރVM�7�	�	�K)���L�$���2os?�d���ҵ�Կ�u]=2{�l�gM	$?�f�;3!=�pU��%M�s�S�HI5~���c>��LR] ʴfZ(MՂ�~�n��ш��&�{7��-&�`L���������E��-xji򸁠�j�+;�h�cI������p�E��+G{ڛ�k��{͗b,�r�-��)kuen����CLO��q:�u	y7�f[�) K���Gg�Gq���WV)��m܀8E�JH��Ӛ��"�&\A������[rJ\ ��悷�AS��嗭'-`*]�c*�O%%��d�?�t�Y��(����jPHH�w��#"'ٰҨ9�A��.+ ��i$1��f��f��EҌV�7�<w��O��WM��eggOMM}��u�7(����.�k|r��\���M��� �@��5�%d�F"1¼:����N�����\&�gܡJ�Q���ܷ~�ME-��k�Ef�@x��H���Fw#2�R|�n ��)�IJjqmmVz:W�L��O�пPO�ɚ�m���=w�VM��4�F��e�1[���dG=y�&T�ػ��B��>��؁@���*@�sl*��`ZԴS&��dP������$ga2R�f#ޝD���2i���y텋��dO����9K�����B�n��*w���cZEP da��:m�x�k�k�P1ٺ��OP��d[�Ѧ�)��hB�b�S^EyA���[wx��tc0���-Ҩ��I��<��"��,�>̽�� ��ա̞�i����:���W���e��[v�_n_�4�Ư�V�?��Q�HH��㻜�z�Ry��""�9���ÔLax�O���a�����!�S�SN�������򐸔T�Ϗ�sp��rʮ����}���+�=��v�0����=�pU��?�
!�ѵ*6@"�NKN�{��Ϟ�ۥ���	��D0-�ߖ"꾁>����1�.U�ý�S���2���yLZ�z�S��$�7e��z�B/��=7}Me���D���:���r@���~(?4?�-�&מѣ?�k�z�;��<���yZ�Ĝ��l[��Z!ƃ`K��N۪��*�������s�/�bd���r:tK���^ōw�뗮�秂Е�6��Q�Ǖ�-����a�����,�����
�`�!�OW����+:9�C[�[���T&���@g�F>�gw:�aok�W�ف��S���OHv�g��MS_; �al��}|����1n��8�>�H�fMJJ��ˈ<��z���s&�7�{���(i_,P.\��
��1�G���~��x�b�h���p(��Z��^a2g�K�yO��B�v�\tS�ʕG���c:U5��W !J�@�tuD�\K�����+/E"�c%�<�d�+h�����;�������^T~�VrF1"A�������|����b�!�~�>]�C1ۧ��_}��߄oFw���m�ay���M_}fx����E�,��?��3�+���r�<���pCZ"b�����RP_1��j���w�=�g����7��7xm��jh,��+#�±�;���޼�����{N"d�;��|���^CCekk���J����Ѝ��J�PM���#joY�ǲgNn&z@ʣ����d��`�
� �<=�4T�W�������������Z�������'ϣ�Ȣæ��حo*T���^�X���e�"tycu�zEA�<u!B�>ǲ݁�~g����'�5����"ޗ�>���oè-����4�e_�洍��[MEb�0����
Z�'��׵Z#����7��ΊA7�Ӌw���l�b�W�g/�m�)X����,8p�һ�|%L��R��{�������`���[�e?^m�=���9&�8J���8�݁��),Eʩ���}653ۡ�Hb�Ҹ�X�}�|�橡����'�3��Kd�0=�����c�!��]�y�i&A�{�����J0�)y�\9�ub�!�N��:�Os��ϸ�F)���I)2>_g�g^-�l�$�����u�%w6����]�ӫ�Z��=""bus����R�9p���'�	N�v���B4�D"0�궶��%������s������,�(r���kȄ�&`�mO�p���hu�P�?��W�}�n++R��qU�f9�mXN#N�A�ua&��H+�^U���P&k��[:�C�C�� w�4__;,<�|{��RA~�Hx������M��i��-�[����7�BEc���:��i�込f����x!����')� 7��OZ*��Q�oK(i���wt���������xx���?|�
H������6☼<f
��0j^M���z�Mw�������0Ѹ�߉x��@?��8�D>�mG/��G��/1���}�cZ"L�(�p��N��@�Ȭ_O_܉�S��DFipٲ� Jf��[�/h"H�Iߴ܄�#�{'�m%��6�4�{����RFF�-��N�н�p~/�����7h����(^��.�+�OG�~���K�z>7L��B��<W���ڤO��$0}�A�ŏ+5/���9,AyA�F|j,WUD����`|8%����%���"�������-�������gb�����wH�c��[��ˉ{��okc��`���Pj'�u��[-��5%V��@�xv/�Y�?�C�p��<Od	���H����N/Ul�YH�#nh ���sDϙ�3 :�L�U U��{1�NN*]ñ8K��uV<Mx_J�Y/ #(�<`uT����z��"�	�	-a�35{�F��2Ϋlѱ5���y���+��܅��u��^����|pZc}>)����UG�P��n �Iӷ�o�|�EI{^�I����"W��BD)A�c��JO ?02s)�[¸��WI��P�K��w��a��է�N6�Ƙ���	[����+W�٧�I��d�{�J�b�ߋ�p�V���+Oo����Ĝ��<�������yq�w:�c!�_���/?��.�fd-�]��^���T�����ל�*r���_N=������kU.���y���AB)����K9���=�2?�N1'>L'4'��Du�6#�hMa�i��CE����_���]@�^�ZY�O��	 �8��<�^;�1��m����"�b�w�D��wL�J,����A���~W��_`�ĺI��s�4=mۗ�!F��N 2�@����+N��`EP��a��bD�z�>D����a$C^|��|mh8���p�i��=:*�u������E��\D��a8�I
�����������E�$��#�����^xq����\�aMT�=��:1a�D��I	�fo��� EՆ5���\�ђ�_c��&�j$�5z_t�Ϲ`Lz��k����E\��}!�re�l*�Y� E�m��v1n�)��$�j�D_�c�3�q����l��h2G�кp����_���X<��}dG�DI),,<{�B�4K�R��M��F���RP�6���@��W��X\�Ҭ�V�b �/Z4����G����]�NN_\**�0�Fzb�p�mږ?I���9���.�~�B���᪘������a�j�mN��fw)�[
���H�
�3U4�3��z�1�u��|��-)�&��}n졪�`FX�e��mY(�;��ŧ}A�B���6,9ӻ�����t��dDw5k��4Q6�_��?��읜L���vnnQ!�/�Eȷ����`!<�'����7C�7B��ⅷ�ӇE���I������W'��LP0_�����	�d�vL39i!��K�&�	5�{\����!-@2)<�z�%.Zy�?�9�|�tK�S6SY����]Q�s]J�ږV#>DY����8���e�mDUX��G���4k���q筓��n�2^GY�Q��|��	4Vk���bO{����Ɔ��:�W�Fʉ�F=�;~�f̗��'ې����<�lε�9ox�j��|:;y�?&}5B��-�Q6�A!6cU���خm�>�)���HM����W {C�6?�s��E��u���s�`}-��o��o5{3�P��	���siX]��sI����������[����0�/���l7�4Af H6*&6�RĐ���m�)�F(�5��i0��Tt-���n��_�K���ۦ:��q�٢�9[P" wO��?kVA�4��.��gFG����Y,�=s��7���٧�wr̭���C� Z@FH^��#�{ʋ/)�����	pDu	����g�ʸ���?��bg��l�Ҭ9��IIu�Ͳ�,�uTqj�>o��E8aMm��/�)KZa�6�Wzz&Q�*��ӟ]�A��I ������/Rh� fO3==,K���gv��3dO4���Ds���stl�[���K^^>����HK��T��3bGM�!/�n�O���7x��k[���jB�{� � �[+/(��dm�"������^m�� A93F�6��y�2���� �Q�M�����}�s�uYU���F��̋��jjVov��?8<�~��QY&���eQS_���K�iʻ@N��Lh��5�ɀ5���x�WkJ/pGh"�m����})#����f��D�@��==N�	p���!2�re�@��Ead|��֬9 p�����h>�1�N4	ڪ�$�{��<~N_QV���w@�������PVQ!��`D$$����h�̲0y��s�lp}>m�A i�+�J�k�­����A�U}O*�1^ᾳڪ�����ej�.Nߵ�OY���o�m%��x,5Lzk��&��Ґ*��m�BH�)�����2��i�P�����Q�N��#3»&ܩ��'�}Ku��pل�q��o���4X]66!��?�&��{z��7��V
L1|����j��*����eck����.�����U���xa��,��.)+�4��|Az�;ʢ��QA_�7�Ay����nک���q��ӛ�:�$
�'�3>�;M��+ن�S~�tO��Y'�P_8�cb���M���+��mĲ��M���#++�1̞0���aM^����4inw����2Ꞟ�ϊX<�B ��֡!^Fƪ�YW��g��K��'��+l4,�l悸Ώ�ȟG�@J�{a����S�?L�N�������z1��a�/>� 5���`�O3G�=r'/qI�?��T�"�%Ֆ;.�Ol���]�c�1����[O���o�OX��a�ņ��t�9���	��
/�<M�EPh����|�h�vK�v��7�"���`z�qu_a���n(`�ܮO��P����$�{r���$�EB�-H$!5/����8�<�RIbw]l���W�!pCȲY�0����r���DU5�KHV6rp$�;2�y�Ƣ��G	_8�Ж{��ۏ"�:ffҌ%��9��D�b�	��V��KC�m��	%"���\?�7�z*��?�3��'TC3C�+���z]]]��<
Z�X
������5'��z!v�]��}ׂGJ!�tx�P��QH$c�Y}p�G�.�u��p8z���
�])���v��ŇE��EVٜx�ˣ=��������9 _#)Bg��X�/�I�����솪�z7$����*�Vy��컭T4��g���D�f�:0`��欫x��fk�d�!�d����M��FHţC������10���˨�� ���;ମ�6ip	yǣ��I9l���j��^��������n�U�Gzr��m��=�b��Nq�^6ǿX2��b������Y��}i��=���j���Q�NX8���S�b=\ay���]W�Q����LA4�RX�w޼K��01�4���9���H*�]hP�����V����u����/�w�Y:M<�����`�mR9%�$�%�T}<j<F7ˁ@nXq}$��H�v4_��D���`N����S��O�o�J�/�w�/(��������z�泚vY��O���ELml���}��S*�ڂ�0����b0��D[�ی����k4������6YT寍M�?�
y�8֎"XG�3
�v�䊭�be�o��#I�EE�84p}ym��P���h�,{���U��W��?��v0��(mU.J=�B��^���;����QdǑ�^��uï$�L��[?�[���k�d�����>���933��oYz*�k��C�ފ�|k%�Q��5!��B` ���G�[O���mTG
KJ"߈�� %��5�o4�N@겞&��S�j���н(�#�6���={��x��vczz���d�̬@U�{з7�
,��J��5�ֆS���L�ӻ '���9���_f���N>��1��Wؘ�@[��}�P�x�G�BBB�#k[���Ҿ	#%#�����h�����6N^^��Q��=��"�6�Yu�֖�x��n*ҁ;&)b���i�Ġ%J��ܣ�+��Dw]b5���F�����9G1��f&�.p�g�µ2�-�I%�>�����b�Á,�k�43WW@��~��/����A�5���e�|"D<������j�`��@*-�Db:X���D��;����]�m����}OJ\�j@5{g��j�M��L{AIɷ\I\����L	���l����5k9��U�sS�?~�3�-'Jro�OWT�2B�;�CA�D�b͏���w
e�Fr�!�/�oՑ����& f�����1�DM��r^�Q���>�~�q�6���#� �)~K:0��o�D+��������5�\���g+��`襙ƙ����J��))λ<)���S�+Y�⮡&��7��4�w��n/]J���+j���h��1=,92CSZ�W�Tx ,����gv�yx&�G��*f�v� �{z���x"�]��bs6�}�Be�O�wY�m�����F5v��.[�L�V��9ŭA�<"m�j�c���%�ŷFJ˔�Y-��fG����B�$�{��U�UX{x�D��[���>��%�a~��W}��O�I��܏�w9Xf�'s��~��WL�Y����9�h�����"}��z�u��F���0��nz��3�/�q���e�ܣ'�35��N���:x���w�.o�!�a�_�`c���MC��7#*�F�94ް�nlZ����1�1����dbJJJTz��F����X��D�ZiQ\���Aϓ�_안�g7��������}�6���0x�g-����,�=���H1P0a����*�H�MibͧjU�X�i4u�3v��/ipظğ5v�k�)�����r��;'�m�<�6���H���Z{rv�6WRB��[���=<(Pu���s��>���^��t�\��۝ܞVU�[{Iz�x�����=B},0��%���
���c�����>G&�	7��(��-YJ�Zw�a1mi��J�°�cje���i�4�B���]0xq7#'8{��Z_l���⣓�*�)�jx��r�l�⮣�Y��A����ZRb;1��ұ;�O��.��cz�����Y[٭d�&,,�/.�F�/��4�Ԟ�`��r�O��\��e���s�y��<ߛt�I:11���LE+�k~')�Y+cz�c��bF�7��JK��R�9}�ְaO��"�5J�E�����2^S�%Gt��E�O"����܊�@����&/����y�
��Z�15ӆ����� ��"�59�D�޲��~���j�2n<?��墲�q�Lf^q軄��'����ʙ�� n��S�������Bo�x���>���?��vp�fcƼ��#��NWRʓ��Sg�Z˝W�Ȟ���Ƿ�r�ܵ��S�5���!y�F�s��̥�fLNx���e?!p�ć�y,w���ȁ�����߂K";�K������ѡF�3���ו'Q����&�wI-sh�k��䤑�-A0��}
'�	ǦYW�鬬���Ppu�����I��� R�NG>���BWN����=>|���݁� (+����>ߍ98֘m�HO�A�r��#��^lmk_��c�V9M�eї���~����/xG�eG�e���bLj#קr���A8]A�b�e?�k������9v�·�ٺx��*Tut�-Q���#?�V�O��S� �·��L��<U�,�L����}�����VO����bo*��P���b�U����!��̫oǧ΃$�|�`D����5�kw�sÍn�m?�a���u��{Ⱥ���U	��*�G���|���Ԛ�T���<2�a��|���[�jd�����R�G4%|��y��q���E�Q�������\	V�P1�=�x�J��+-�` 7��&�Q�h�E�dN&}nfh�=4�da�W�Cų��~'V��}|�-�SRt|����6	�}�4Ѩ	/���E�퉢JUn�_�)�tl���<�"��|Uu#cH���6zD�/:����6���Z%�_0)C.VnxH�^G$��#���l���"_h�ΖQ��'5����۬hzu�s�,j1^qA��s�ض�,{�+���;�GR�!|�9k��fF���G�G���/�r�w�s�@,'���e�],�wf�j�6�#�_ٓ`�"Cv�K������g�o���,x�42E5@B�kqh~I�3�JOR��L������<�����G�x5�5к]���4.��,��r�AN�X2���nFtm�D����tt����
j�!b@H�ezs�#j�'��^��nn�O�Z?�M�]�j7|�~�lM(�4�N)�&<|V�˘��������1Y�j^,�3S᱇�Ω�5���Ix���c��m�C��Y���PG�s���%7�����)Tl�cu�K��"*��)��hQ`���]��R�r�+�SMT��mk�5Z��m:}�D���)hZOO�J0����-;YY�*{����S�%-T��,--O.�lg�����3j ؄pfvv6�E!��^W��!&Ʊ2��D�e\^�+�V�����W�v�3�j'�b.����2��17MO���qF��Ȩm�P��P�9�Es��t�μnT�s��h��&ȿթɸa4�##�ɰ�WG:V���E�u��T���w��u�$+PՉ2�@ �LT#{{nG t$ɣ��oT��J��;�
��~f��!}����ENE��� ��p�����@#]��<Ώ��(�r���l)��)���������3m2QE�qR)m��Je��ys=^�	c8�H�q����ޕ�	`̝X3�ɧ|!���5K���XV�,�iE�����������G�+'R�|���iD�h��j��� � �ڢ{�:��w)�2�6�A�?4?6�n�l>VYݛ��	L���L�����Л���^�bF0	
8�B�r��So7XЄY����~�!/�#����r��{N�����������	����@�G���ޠd�8��G:�&ga�;bf�9���F�����JjA�s|��]z
�\o�5��6�W*����&��O���]ܛ�X�;Pmu����I�Km}ј���@�W
DB������nE0lu�x��MО��^��ʿ:|4O��+j��֔�7���Aˀ����炢��. ��6�����ۊI�3��20DSڇ�����K�g&�®S�v�J�pIH]��~�4 �:�|V���	?O�$����N�����4�W�ݧ=�s9��������|��m�sZn(uou7���jpl������9�KZ^�\��5N@��
N�e��)��߼q%�#�U���g`�t�U8e4�-�l�" ����������(ӵ�����p������䤈�o��+��Y����.��r%)[;sRva(L���Jb�M�qL#/�Pa����	)��l�ow7bW�p�|5�h\�Ul�r@��= H��V3AA�vzz���l�Ȟ��-Tq��N0�A�'������Zy��g�J�mD�i�ޔ�4�]]%N@�O�	��k�
o��A���443����y����i��.�(Ս���踻������t\��\���|ki���^1�����VQe�Kf�XX�~���>>~���E%�>�0��؟�*u�ݓ��J��;���g����/V�Q'"��.cPj�مB�v G�!�;fRd�j�)�r�V�FpgH�Nd�e A,����w��M�ZI�_s�Y�hh�9�s�z蜾�Fpv�'��=/teM��&���a����M۳�A˶��k]-�e�%��/�]�/��;��ߔNZ�e�.U��O0�3Ӿd����y�8�b'����/�3	D���V�c��!���o>�~?�1Ͽ>B��u���e����]m�N��\V�_z{�{7�L3���O�ܑ\� *O(�5(������ݜ��ʷ ���R$�<���z���8�},$#�Y���|�ɋ>�㼖�?f`� 0�]��	*�*&��:M�au���;��n�lw�ߓ�=duy�Ί�3D����郹���&�w�("?�NΈ��� ����5h���b
��ϛ��L}l2��콲��Oe��.�n���M��QQ�0q��&_ُ�a���V��s�aQ3��>�о��P�����E�������~��.���3N���[߻��	����9�:Aۉk�����)�)ܛ�}٫�_��
^��u<����N��KI��)������kw��a~c��N2>���$��1O�x���W1��#�*rқ��+��U	�c0��-��+!�c��
x���� 3��ۊ�Q�����~�]�p�����R~w�B����Ү�֠? ����ySW�q|�w E_ڜ�F@�B;G�B�����"�g��=K�>�Y��u@V�<E_2�ES���X��gS�[����M/����W�ű��F������b����Ql�qq<���f|�m�t�x�3�1��x�ӱ�GZ����*��ۢ7E�49!�^��������Sz��٨�<Nڸj�D���bC?J�� ��ʿ��͙��_�bҖ�T���I"�Õ�*�� �����V��.dP`��t��l����e�7�%�����nsRR1��I�?�=�˄M����mLAܟ��}(((�w~#���.mK�h������p��ӋdeY���	e�)U��=�����yN��ޜ-E�>������Hǒ������-G�ک��S�/.���G����H�s�4z�v21LV�e9�[�9s�fX<�u����)�wb+�3M�C�~��?�~�wn����8�:{ؼ��!�X�hYL�r�O貓/!���¹�8FZjIl�c��d����Z�\�i�2"�Qгf������sJ3��042�g����C�u0E��7�
���7�Ө���%I��O�I�Ø.>�r�mX`�g67Sk��]A�k��'��1�2z ,26[�gr�v�붵S�a�7��f���G�?��#nܴB�1^9��"�l�&���f�L6Kd÷��q�~�~���Y�b'����l���g��`�e�d�����jM:8;kPVe����}Z���R���X�9��+����uduж�˖��+Kb�c��p�*�dE�_� ���D��fP�*��B�zX	�D����(��ʞ����[�M�$E��U��q˫��۔s�Jy��aU�_%���+uj�9�i����A���)M��=ßk��W�|��s'�Ѷ�PN+=c�7�|4��z����~Q,���m�ǻ5ɕJ��&wJ��(ݮ�Q���FC]Xi�$#;;�	���U��;P��-Q������5K4�����~�k�x9�WM]��p���C�6i�f�I�t�ĿCD�/э�����}k�{(�}���au��ݼKu���9	�M��.��<���U��0W�;Ӻ��%�޼	��>Q|u��X�:7[�B������C�T?�V�j:�z;w|�e�\��\���7��[���Cf5>�X吸�ܯJ��m����H�%�@�"�>��?<]T���QZ�$���0&���tII����t	Ȁ�5�T�0`�QR�kt�?���s�΁���'�{������k���lv�e����@lc�s;�����ǐ�a���IBF<'&J�+�W�����PmM����-���UP�ku�/z��YO�W��Q�h��U����ͽ
�e���q�1 8v@�n"�ے��m2�����8�c��5�8�9�"��{?
����ǻ�1_����zᵬ�������/FL��K���6�~7@��|:��em��tO��-X���f�Pr�7G;S��퓈�Bږ��c�ݸ�˽,~zÃ#�W<�'H��΄LO����*�D�x�*2����76H*�^�鋖���ZF9.����g���JL2�PE����[.�����*"[[1���Z��\�m��0�|���w�/dT���T�`(O��k#�y���;C2Q�E�Г���V�� )_�Ol_��~>�jm��	�)��'��̻I{���F�-�h�jœ����ͨ�{%S�;۫���e��5�R��}����:Wm�T��Ԫ���յ;����xh9��[���.��eA��=ge��|�F���J���t�x�idYA�*��F�Usdx��m�D�^��E Q��BG�O�ɲ6���h�n>:1d���7l�����ʎ����D��"^.��8��Ţ�o�ͺ����ge��S���z��w��?�q�"�I�w���ޑ
������j�ٸ��r��䈼'�Y�B:�>��b�a[7�Z��2�.�3�]y�l[����+�;�V��oF'�.�������_�����fq_�G.��7�&�^�΍S�#�Yd=FFF�`L���<��:I�}��浨ʨ�8�/&�w�"+wG�U��P�t-Io�G!E�z��ezz����dH��e�ע����7�/6W?�:�����b�Ig#�>�D.J�}ת_�����]���H���t�iBRLl�����cٱ��$���v��}NN�?�P�>q��o�kr��{W�Փ�2�+ج;�IQ�� w^+�M�{��?t���js�W�a賈��5��_��d��ܑd��~."�n��x��*+�Fc��Ÿ]��Wv�8:�z�<*�YY���ϥR٨����7�E:�=��������_��A�V��rZ��y��(977���z1����������-oD*uӭ��V���t�EEE>?����c�tuѕ[X�����_k�,���2[����%�dC	*����x���awK-�?�����1���+P;��'��.!q�g��y]GX����1�By��[�ÿ����.u:�w�7��b4G��;)n�(����srjW%gfaIW����Ժ:����U��'���׿[�;R��2Lgu[����S�E(�^&{!���;���nK�ŷ�����v�k��'���Yd�?_f�h���%MCq}����2/e��� 22�v؋����6�
���u�ZSĩT�`���x<K�ƍ��QԥԴ��~9k��J�; =^�w���pX
2�J�W����Û�|J�5�jB��)*|��Wn@SҮ�H�[-C�d^�0~/*"��4ےq�DE]N�fA�OPq+,
��xl�x8A�9�fs8���1�0����G"����ӝci���aM��~�u*��͘����i��Y���̫z_��j��7̛���l!�ڊ��ޞePPQ͹�֦t����c���
T�턥D�WLlik�@�1�S�n����3��Ϧibw�7�<i�C˛��vv���@�C�f�����w�Uބ���ׄ'|u|k>�����7�i��@]C�)���'�Fv�L�����kT6|��X���ɺ���rl��������e�,--�d/�g�$N)^��;�l��T���e��
��s�Gd�-.Z1����뱙~�7ߊ����٠ܤ��kJ*�1{�cEN�t���VS bߎ�Է�M�UCvfN����$��RT��L�ǧ<��+!�b�j����f�Ʃ�4�Vwb����!����,�)"�u*iV���W�H�H�$�]]�2�w_������#O�LP���uuu�Q����9ڻ�jٵl��Vy�bd?���.^�ݳ�h2abbڵw�Sɥ�"۱RR�|�<H��}��O�����K��߇l=7&j� @�������MGB����_�b�:��^m*�J�(�Y��JO�)Z�v��"ň�E�L� O�K�Q����jge�iւ��J`Za��k�[/�)��n}��}�����!��䣏�f{��;6�ELy�/9��#��=�j�[\\t�t�f�$�q��p ��da1�<|���� �u����#rqY&�Zy|/���]q�л��y��A���E�Ԥ�2[	�&�>�~�K0[�ǏϠ\X=<D�ۚ�bN ΓYJ���Qϑ7ƽ%���>Y����ŷ�7ƭ���/xUE�͗�i����Z��3���Y^ޛ�/+�YY��b��*Y�Զ���2b���H���Ze�>�R �x`����l�1���&*�L��''�"bb�0�TtB�3V���?��w���\q�mG�3~�����&0r�h��gb���KI7qz#�N��;S��#�'4�覐 R�{�{C���Ij��f�?�ç�@�����1xベ�΄�!uh� Q�C��)�FF���q8H����yS�|k���D@:"�k��R��-F��ի����?y>f4r��zLA����sHFvY���I��i���Ej$�uE�i�	�����������#��IT�}��t����#���3���.T�N���U1����'���sa���_R"�m6,V2;�trsҳ=z�y��؈]{TSs�<�X��0�s��&?T�s�5�8b	TO�����8m�N� c$d1��fT�H+�>ST�����o�5C#�5��ӽ�B��'�
ǜڐ}]
�D�y�e6͐XJff����4B�J�6xƛ��JO����-͸=45�lk�'*z�`}��ug��wi�4�����8m�D�l������-�T�^b��Y�鲌{'&c*�	GCin�ż�>=ԶO��ffR(�6�"&�uQ�z�A����`ڴ��a�-H�5���Ȇ�����LaϯW�6��n�5��/�|��34�|/�j`d���}Y9D`�f������~���f\I0+�Ϗ�/ʨ4��"��F^�m��D�����=�FQ�I���1�T�ȥq
@�픩Ƭ�	x9��nyIpwk���!*�����:��gE���6�@�J�J!�x7����%<d��N��,��D"6<��K)����z
�mV���@��:%$fߑ��0vT��:�<�4/>�t���x41�)()�������`X��Jn����F��<O���ۯle�Cft�7����RӜˣS�i��D�!�3ƕ
��lX�XUQ|��V!-��ѷ��4�$�\z���/B̍����3B�p�-,��K�W>�N�8��1lhѾ���;H�%����Н������v�w3�|�X�k,"���l#����p1��Ǒo�.�ۙ��t�>]�Xm }q>|�餱D�0�%����&Ux����>�KW����|�������w�&=�����5�����ΠUt"k
����B�ʼ,��6���3�)k��q>�P��Gg"Uc�fG��6�A��#�6�,�C�{T?�sƿj���1�({��巏Ϲ���ݹ�Ԣ���	P�Ξ�!_�|��X�x?ո��`��T{R�u�Y獎�u�2�K��q�'���?�+4��B{�����qi�+���ȱ/9�S��7tj]�� tN�;n_�� �(I�+VZ�#��\"�E�/����tec���յc>/��\دV�ޣ��f������&k 2v�rh�(~O]�RD���u7�B�h6��$-��G�x���'�8K=��~`a�X,��=Y%�S�#z���ř���U�x����7O��m�;_�[_
���ux>%��i��L��]�]I � ���_����C���1�i��p��i_��'�TY��B�k��c1�k��Wrl6vvv��6U��!�����)���CL�*wE�y�|�������padcʮ-ch�O?�{s��J������w����O�#�Jx���+>�}֡e������Exiv6]���|�5���Ёl>;):Y�U=�y|6}�8Q���x*���c��6�|984�Sئ�q1��W$���z�D�����@U�KqC�8�h"r1[n����[�M�<�gu�ͧ3.|W��2J��} ��dM�\ ���_��HN@��K]{��������<N�	W�ܖ��9���d�� h��Ε)��/:��N-������Б��[�8=�������5�Ą)?�ri�{�"v�#��zH��"�m����c��h֫��&�sv���j�"���bt�rm-J����S%[=)ny�?����A���3;�k�i�������V��w�$c_�~Q����۝-Đz�:��}��Y�	ӋW�\�W��M��K�ގA��eq���i�jw��ܬ�I���g2r�h0��J���(@�`c�y�OC���.��9[���,�L� beg�d��ڐ�j��B��W�G�=׋��D�|Nx�;�4&��F`�Y-:1 @��ER�D��fI�K������WQݨ�Z���;������%LK{����޲`H��\�K����X�������F������
tz�ˬ|���'�n�F�7�����98z�L�܎�m���8�%0�$STS�_��ʫq՜�A���J��5�(놫@L#�+��e���&�<��5�x(.Z�~��"!�-�b`�ᡷ�x�U}җVs��5#�9����/�?եg�龙J���g1��Q��Fƀ��\
��)�<�C�E���?�>�.H�.�v�E0r�Ȁ��`oD�ƈ�#�{��<<G�t�M�Z�w	��3��u�~B�+K���vgބ�ff+sVo-�
%�ޏ�{�����<r`�F��
�#��`��Q9�j���v?�]��Hv�k\^���*�����}�,�#��i�h(��<�{쫔 �쯂ʦu�e�d&�c�q[��U��Fw�?�E��Q�#��X:��Xȹ���<'Ŀ[���0�����]����NL���J�_+�afN���yS��Dp\ׯ�Q�!)F.�O�0�e���aq�|O�,�u�,���e���iC �a�'�(��%:=��2# ��m��S����de4�ݧ56�>#�[����(�o��V��i���@r���;ㆪ��s�0�L�鼜BA�i��+RɉAV���V�RTT����q��4��V�d��mm�gh�1ׂX��+�vJ�0�r��7*���4���u ��d��W��e7a��l�h��m`͚�Õ��-��3v���y��	Ǔc����?�2����:�[�|x�6?8�u�{[����XhHI���2�N���!0Ž��
�D9Ԋ�|��=�(<�d @�dK��LIY��$6�b0�l�v���S���!a���7�������A/!i�B8�u��I���V�~ώ��y2��f�w�5.��n�Yb�`����B�8�x�j�����z�tY�`�X�g�l�A�j;�M��:��Ɠ5Ԉ�g�x��??�3�{�6Ɯ��/�����hx���O!}�4i1ז�-F��L���A?��&� ���?o��L.�_-��	������=��W�τ��iC.��
6�u����W�����}A��i���2�!4b�q�f65�,�R6��iz���K(����ee���:����7�P��ı׀>�o�`�,�����I���,��%%W(�m�k,�y����0�mŻ�����* K�G���Յ��!{?�@oZ�w�|ʁ�on�v�� ∌d�`Q�7���@qQ��ٳ�n_�Wd*��;	2�ɱ%�4�B��]1`�,'���c����55�W����Eߍ��x�?�!:�����.����r;������ѯE<�u>�I��םPt��Y荐e<���Ҵ�|��'�|,���T���ܱ���K�m`���YuD�*@E��dO5�^\EG'f��%������ Ntp��I�o�����>�߇�Fu������3w�d�T%}�`�O��:��)�h����1.�Q7�o��A�8- ���3{lL��C��֭FE^x|�HK�{v���9uF�8Y(s|2�11]��D��h'=��)��߹���ʺW�Ҽ���	�UN���YVAթg�gy�j{j\��&���ݯ�\��V[��|��j=>��cI�}M��x�u�c��Tr��Io��^���}�@�>�|h1z`Zm����۩��BYC���\��r_"���>��<�Kx�L&��J����e����kmU5��T��C&qAq���1FsN2z�-���J;�u�����W�߇{��U�6�ֶ���y�\;�t>l�Z��1���vk��X�:_�j�M*+"�3)��Km+��@�������"����Z\' u�����s+dV�I+S#}Fu�-����%:Ǹ�	� &�?�Nʔ���kV���>�w����ET<x� L;;Æ�o�[
���o1� Y��$yl�8����$I�5�* g�G���ZN��(n�1O@^N����O��0�5�2���+���ᕡ�&6��oK]��W�\a=����Ҙq笵_-בt��^�y��e!61�5L�*�����~_O�y�ym3�n�`�������M���ȵ�K�ѹO��6�����n�-=��k���$��ͤ"q��Ƹ������L]v; (�+��GY��'*ӣJ��0��T"Yz!,-���?�ͨ�ݟ�EAx�R7%Hu���ݷ����f�+�����I-��c����i����T�/]�y�FD��6��[~m-�i!weX�<�ꚫWIh���<藱��ͪ��Qʤ,�R�֫qtpE���XrR���������@Ha~X/��� �M��}���ߗjj���e��M3@�,onr%�$�����>�%�GGGg�[��5��H�n؋ܼ��ۏ�2�w�< Paq����F�ZY���W�����9����"^rr�U뚹�L���o�(y�7�mR2Ň�a��bbW���kO�C""~x:C�G hj�R�<�a�ܼ�	a�$R�Om)8�D�X�$�,�D���=P���7&kH<� �A���e�h!oU��%]6qO��Ƒ��%���p���5��e^Gt7�⇄ �(I�z�GC��gCj�r���=>H|��"8�{,���t��ú�>��PD���i���{�@��5A�����h�>�n�X��3�=u� It�����'�&���u<�G'1Z�)�X��#�1�����^}�	�rbmmqj�E�b?�ϗq/�Ǽײ눌5�kk˺�R�t����=�]��L���zr���j�uN	��ڈ���Ku�l7�7mRNx�h��(t���~�2�
��8Y0�_½�!�?��v���x}�S��i��_�3z���?�̻�HZ�������L5s]��Y�=D���F=�٪1[Z[���~�Y�b�Ur{�}�*�}HX$E�M���LKk�/�y� +W�A_u�΃�p�䫭�w�4���ϔ�N=�@]�Ώ�(˙��!W��0��T;���  �T��|�
���YҢOEDBb�k�HU��ʬ�b�����U�T&�T|*��W��n��g3m ���n,��!�v�S^fƩO5�nx�i� 9����}�}�`z���[��c7K�g��f��Z��	��k���t'<�T3@����;�֥?��ʱeJE�`�,�CBC]Vd�b����x����t�����>�<�ث}�^�Q���UdF���qf����7�����#:B4.Y��i��.�h
E���$i��[������}O�T:Д$�~*����`$����k=2d����n��!$AM�.�W��.,��o��c]����l�)#HK����0�����l?t��#���R-���q_e��{�n��N�@x�E�{�Sa�;]j��V����G����g���,���Ԕ�
�����M�
!=�&fP�G��:.���Ϟ��e[�19J����4�If{�0��64�Nx���7'x�Q)q�s�?�dPX>�tB	^	"ZqOm϶7�=�݄�O��}������f�b����9�_뮎��lnnfƏ-/�\J���n��ط?��5o�7�j�d��r���K6{X���=�v��\8<}�l���oC?����ϕ�\��*�?�l�$6C�U�Cy޷e�̱&��ZW�i���#rg	-,|�B���Ŷƞ  9���n��0VU��5�4��UfS6/��4�}j�6��e�h�v_bt~*��yx�M����s�XSB���G٦~�%\]��FB!+&:��p�/>��Ĺ�j0;������"c��f��⠤�{��7�j�x]^^�ź$߫�^>�M�V@ZID���x��=�32�-@YchH��H؍D��n*�
0i�f'Cqs���[0�:��]~�OP�O�����'i�C�!AV���ÎN=���V�0dI�;�����2�b����Ⱳ2ڷ.�G��J�l��u|g��)�����։�����v������s��X@������ۂ�cqK�\�5�3����T�
/�me5��
�Ӓ����I�ϡ��`de�l������ߢΥSt��D*
������Ԉ��r�0腥��亂���X�N�|޷�p�݀�tvЧ~-���U��m�l�,��E�wY���+���Ā?7<sm�B���� ��و� I�_��P�zd3c~��(5���#p0TP�s�m�2�na#K����!�`���玷��o��������~�_��z}H�Ų6p:�Y�d��c��1�ŝ;DRЮų���;̌����=��?(��UU�߹s�׼���t��Af�� �+!���d���m��D����l��吝Y�#��3���g,���������5�B��0����KIߒJd%�敕ż���^[�PNIO_�L)ˮ��2H?TH��	��M%�*��/y����vJ��͐���.ׯ��b����8�,˃`i�̽m�յ�w+?��00�p�"+g90��A��1���~*��4�s4��Z�[o$u*h�eeOfQ�Zےem�WE�KZ8_��I����C��IIS��U�gn��۷ϥ��i�	���3%f#�6�@;��N�ߪ�i�� �hHFO�k{a��-��.~�jB�^�&�c�l�2奢��L�,!���s����[��^��34	�
����}xg2S�[9$���>5&&����Z����X�ёT��1}���~��ͦ5�g��Z����RC�4Q�w�J�����kk������+�� �b~o�¤�w��J��Ve���5i�fӴ����\ֱ�ڛ���>�$�@��^�8o96O�`Eեe��؂w��-�å�mZ����/"*w�G��ܡ �s��j��S�Ⱥ&���O��)1�e��kҒ\
r�\�
��2�>鲯=�8������z.�:[q���w�Y<~��1���TVr�ٻw�/�e~~
�G]{Ƿ��곟��/~ �O�L��<�p3Z��j��i��^����{}L��U�m�Ik``���n�v�! ��$:	!����ƪ�ԇ}�r+�!�����f��&x�iS�G�����{3���i?�y&EK�UX���?:�+:iR�&�5\���,�T�0Hx�mM�x��NY����ge�KXF�3��O�j	o���8���~��~�#`�*�X�{��2�+'�c�06>�T_���܎TRc�K�ߏ���[��a/8$�}���!���,�a3���2�M�ﷲ�ӳ
Ĩ���E��6퍾�����
�+++5h������C��"=	!h}z�սYӡ�O�Z;��Xc�3��uiw���\v)����?ڝDbͶ	I��&�u@y%%Q��Lj2 ~z��R�R���<|[�i�*=_K���Dn�L��:���!uxsj�o���w�k�ScA��7�[������j��B�dɅ�t֯�;Ӂ�B����"Է�R��\��8�������K��`0H
�M5j�jiQ ,����a����
�o����͛���~��"ֶ�A��������R>�Ն�`�x�l�`w׫�2#������&�O,��|�1 Ϳ�	E�#Y�O�m����8��2i����O��y9ݦk�b!%���
?}.�h�\�y'Ȋ�477 �<�'�":��n�>'|�a6��f��>PN�Ks��:�d��Æ�*�k��@H]n�Ϗ��Z}i)��3����mI������&����J���ژ�@�ͬ��[*xۥ�?uS��G?��p�瘘]$� *>� %��Ⱦ��Û)�IJ��HL~�l,/��8BT� �֕����|R\���A�E��({91�*���*W��57O(w6��J�>���}+���6�:Rd�W�C��R$'�w8�2�r�;(����Z��	*0���/	yy��;�4o\�mU�4y�nA𧀲ݞCB\����ћTv��>��c^d{|(R<�J?��G�N���8�r4��r�-1��R��RO���|��ᗼSH=��rI=_w��uU2z����Z�Q#�����Op4�*!��3 n]j�W�����zj*��X)�K{oϮ�0*��-v�fгK�������TOHI��jg#���bn3�:'���٪v�`> �������F̌i�Y�E�sNa�?�8�\\��M� )hKKf�����X�a]Dϧ�������*�b;ۗN����I{!7���^.��8�oir:�Ae.� �MGxQ���'!@����eJv��m>\����n
�n&ݳ��0��7!4���W�f�`�b�n=-��W��~Z�?���w'�|��Dl%A~v����%y�O��9����㑍a���D��L�!JdEl �<�m������:t�[�4mQ55e'@O���x�#C��u�5�e:������a<d�Q��~<4^�JP��!닠~Y�N�5L���_�R_��2D��f���{�����$JK���hJ��S����::r�vS(���yJ�\]��c�& ��3ix`����Ê�؊\%x܂��>l������Az�iԬ�;�1������)4a��m��j�S^���JR,����](!����P�\LhE�r�܊fi�U�r��5Ge�?|�W ��;X��Hq��n���P�Y%����SX��75�t��L*�<� ����N'��GFE��.����}��Ӵ�3�F��%+!?��TS������Q�P��
��n"�D� ͑�	��%��S�d{�s�[��`L���3û�QȮ���HX�O��������g��� ������?I��7����x��n�����m#	Jc�#>>��R������l�/ʟ]�|ݧ>3.��;��^��K4	!^p���4�ֆ�M�Wٸ4NMz.Xg����iS�`�ڴ�����b�!�#+ז���c֥�^���=w�����0B��l�jI�}C@$�]_�,G�N�M���`�iN�!�L+S<�af�ڂ��N�8��{��"n��o�l[�X��6]}?:��r��`��|}�9�Eݡ
����}��g�V
��~�o�qL�fc�}����|*���+���R�Qa�W���B'&&$ �
����?�9��ؚu0�U*w��8E�͞|�in��̭n�vz/J����g�:%���LB1&���-���"��sÛDYZ�p/1�Sk;�ܽ�D���ta�u��^(R��2�T򩳲��%ҠP��U|ΤN���e?P4�
:`qXg�>��]�E�m���?���dd�6���z���4߽{�eʭB�J�'�޼���[��`�D������Ҩ�����j/�T���ܧ�I��>��a�Z0Zs+��8��?MMN���\HNy�|�Sk2���8�����Pq�d����Y���ֽ�:Y�^�v�r.�W���Ng�=N��T=|J�|6��Pr���(S2݋�+�?��㴯]��f��	/�)�A�E�+F#9ֽ��Gd�(�,�x��`��r����ܜj$`��)�֧LG���f����n�Q��~�X����J�4R*����X�������\MG���
;[:b�J���]�y�bT��69��}���ݎ������47����DΞ��RHw�{���#��Zhh���jQ�S�J
����٩p��)dj���zP�r��kaP1��zLj�h&|WHY�Z��������-Q�׿K@��11U6��ܨ�P9b_�;?��&��*/�s�
���k�0r�liǻ5�9����K�>%��า|���D;�u^vQ8/ݚ�n�d�ƾĬ��7|��Ù�`h��(k1�#t�}��=�����J�4~�,�_ɴAː-	������N��,-�AZ"DN��VR-w�8�Z����l��E{�h��?�@g���>n�-  `(��X�̧��dd!KM��1��_;�h���|m���x�|����2�H���b����PҶ�j���%+��C�W��h�3���(�9���=~e/D�?h�����^09E3V�h�*�Ȱ�V�g��i����ko��^�3������G{�wY�MOO{0;���7m)WW�sx�`0��)�tBBnd�kc�-�.�P��û*���Ӥ�:�%�A��RCrx�=:
�kkQ���fɟ-Y�21-9Ύ�啕����5�c�sI&����'D\�x�jv�]\���m�]>��=Jt'��0�*d�5�d�����HI�z�[ �� $��2�ɹ��x2��
�H�54�j�����t��x
 ��8<��y��{�o���nn�������%%Nep:��\#Vz�j!�zkX�qk2�!}s�0q^ʨ�ټ�"<�a͗����bY���NQt����+��Xص��x�TF�Τ�פ�$QD���Y�f����1�''>Â��="���u�:����4V�1�g:>c�s谸��	��/ol �Z�uw �G�L��N(��C�_�Y�졍��L � q��@X�ם����)��0���&)u2;}m2UŎ�IŤ�9(W9F��{�`�덆��R��l멣3���l+�r�{�P�_T���N�N�3W,,,�=�/��尨x�˂h�Ue+�����o�޺�&"0yP�[{���Lom&56�96��'�s�EPnt�%u�L�Fp��L"����SBе��M���3�O�TB��d>8� DR���f���cG�y�ִ��1-���,>��g>9<��1���9b$��Ƅ�����.��_�a��on:-T�~���pe�<��l�!��)y���Vn8={NN�oh�ӈ(��f�AQ����?H˪�������~� M����;����8}@c5!�?ͦQ�r�8���(���V
S�m�/ic�ȼ�ч�>�G3V����J�9�|�a��b^.�@}�\K��� �p�&s&�|��j�6�]?�yB*������`Y:�Z��&&t�W�R����� �2rr�5H��E�>9�['X���@B��9��Ԛ����[<��2�l����LzM�æ9�[�~��.��̛��Ov�r؀h��U��A�i��v�2o#�O��$� ��s��t?z|�?J\s3�X�V��7 |Y�O���'��:��vrX�+�v�<�_��͡��7=3�*�ʮ��B��݌�-L�qu�`n��X��P(���\NN^>ʜ��̴Q,*��Wk�qUw����!7�G��1fA�G�_�.t}(+9�0�<;A_vC���;F�ؘV�󮻍܉�)i
x�PKS�AG���'�JTɪ�����</L�w<!�llt	P�����U����~��K>=}�Z�"ﶹ��*#~�3{xJ���9�=��ࣤ��=3�\���9tz��I\�>��B[�~��gK�ԼdA~���xu��vj��zT�ozN���?":�[��ݾ�!JEW� ۈ�i0=�`����o���BX��r��-�į�&F�@(��t�
�̦���h-�+cZ%#d�c�zz'������q�y'����23#��f+DAJ��8m�q��m�8殞o!�������KO|_(�Ƃ�@Õ�eTV^�}�Vǻ|iY����F�)�<N���(�^!�Zv/(딉�e[!�>~�!��N����5����5M����L��3Ǵwⴑ��w�:x Y��g��{�n���\�������a���2��~��*!���Z���v)�k�)���}����n9�"J�񀍙'��Gol#�>��!e������\j���?A�F���봚�Z��C$�c�W6�� ��]_�૶�]z_��`�H��k!�؆�j2��~3�~!�ȘD�V�d�8���Y���y����N��M�������昞#�$!ӥ������kW�J&����r|�|���%;�֌9��{K<|�?�=��7�p2=l=@�̚�!�^�6�u�j,.N����ݻ�uv�*��{}�m"��G7YeC����j���ԩ�s����s���R�47��F�8����u���a)��/�v����%�]ea/�i�ᧅ�F�5�"[א�)�т�F'&�*����^P��/*� �|X��������;�0��*���`~<0�q=��&��� k�Gb]�y���$B��H�J-�\�\@6�^��ʭ�6�l�;��Y8�""����M�Iн��]��V9���v��j�����:��Ve^`�W�_�Ԙ e�T[�Ӿz���c��6��n����&�0��Д��G�v�[����=��V���Z*I-x������+4ij�H^�BS�0�V��M���$�4^̄�Ȥ���h	�:��}�V�H<���>nq����+��:J��b%z.tq��vW�j
M�R�(�'�̰�E�v�1n=B��	�>�s$Qlm��]���̭3�4{�D�-��Ƶ+k�����ߚ���h�-w�{=�����\�7�F����ho�@��&{
w����YP��7�(�e��L1��rr8� ꀲ�乌a��{�O/�%%S��o��6�p>{J�.�&J�Ze1&����Ț���{?ٹ�7����w�g̶W�W�NЅ'G]R�)b���Xe���`S�ut`�
6�p�V��c*Ep��Z���zvY�]����Y&t�+`�/�Jh����͢����(njcg޲���O^J�7u�]�W��!��y���KO�y�.Wǡ�ӝ4�p�f�uK&�SS���Z�a�Ay�ؘ������Nn�+��<A�3e=��Gi��n��}��K�d�qZO�(�dkW�b8T���|-�!yu��e?�'.�bVΖ$�'0���|�BLS����ELϿ���As�#�ԯ<�x��$��p?pt���Q� ����L�^�[}�Lb��47$��Y�����e�j��$�u@o��L�s$m1M��������d	9��"��[�B;b^C��g��%<߲��kסC���3�g]Y4�]Y���"��i����m�;��u�y2.1>ޕ!�_8�d�zz�ߔ�F�ş4�{y�JQ`^uM�3�#6Y��u���Fی�O�y�Y����b�mp5-1�vPkCPX�[1q��nm�4+oooPLaQY>�ً�;=W{�w���-U�u�������e�qӶ*��:���6�����		�M���J�[�Ȩ�W	�=�`(��IJğe��؆\�(vY���Ao�	���@�����T�Z@�,���R��O����g��k��<�~S�����K�5i��M��u�����O�O<��y�=����^YY��"XSR#�����/��Sm@�`�֫������9Wu{�a��Ӝu�Sg�C�Z��X��ܦ���!�$+���S�\ 5�m�
�J;��R������}i�]�8�k�"ku�5�=�����O,1m�>dۉ@���I��g�!��c�u�K\B:�Ժ���#"���h� 0�5��(���ڕB�O5ba�����i���JC:��ʚ�Z�ho��l��z+���ڞ%��ᑄL�fM�`�#��+C������?�U�qC���z�,]f��ɱ �9��x2���_��������$��Iƙllz=dde͘�o�Q浒��/�瓴���˫^N�φJ4�-W���1�ϑ[��Y'���mW�NV��e��K��6��x�����R�ϵwc��-q���Z�j��'�FG��[�������F/��z���F�%�1j�,�ٶ�_�����i�n��w�.��T�ʇ��s�tv����W���J,��?��qj?�3<�'CǊ�3��e�{�.J���E���������(��E�����D9k�Lv��~%(��0_��u|�C���AE�=�e���ج���}�W�����l؏}�b�B���V�
(�l�|ؠ�s��u��̜�Ab.Ud�I}j*I�V5\hg|�1���pMSSD�amAQQ.�Gѱ����{���z�z�����I0 :��iVΜ]�[!j>�A�=FE�%v��)u8���ec�̂��6�ɝT=���kl����>��K��R���1���<N�� D��ۊ�}��{��*^���ŝDٯ}7�ӛF� k�b�8	����1+�Q���ak+�c��a.���L|En/cf����t����N�s�������{ÅIAR	AbP	�n�Tiai���E@@@D�A��;G$`�a�!�`h�A�����|9��`�b�g?w\׽���4���܊�H)�D��z\3�ȼ=�U����@5 �G��)(�d:ZH��%<@EMmlT�;�`�����:1�U��8߈=tdqF_l�m�Lm�D#��1ocb��W��%q��5X@�m�,���%�/�}l%7���P1��96�͒�s�_ψ�^_ņ�pDa97#�q��}ݣ�ܜ2�j�����ǻ(��6���<�J�.r��.΍Q���	�k������M.�7>Y���W,X�h"߹׿46��M~����M��˹��4����=6�漶,�m|�/�3Y���E�ܷf�xʧJ� 6^����=�x����s�<<�`����,�vyߖ�n��K���C�
y����L��ȑ��t� ��lFg��dz�[&���iibС򙻘��c���}(��r�}�hm���l��1�2<�e��e����,Z�\�)m�ɬ����Y�������g���3�/���p�֏��F���P���W,ވL/Q���z��,���jE%%�F	A�~b3A&n��\���)i6�����i�l����GZ?5�]_�2��5IHvsss�M�2=#���5ap�WD������n$'��N�$0o]"����~$�{	�,:}z�i˵�|z�"�6��.�8�K�r��X1>�9��^Z`�G���(e*?j]-C�K	C��b��JK�*+��n��[�N������U
�c~!#���.�|ʘ�^/x�ĜI��uyr��Ƙ'+�`ߢ7Nb��y����牬ĢJ���$_f������[ !����u�m	�^�7֙�u��,ӥ�����\���ӹ�ؼ/��}�\s��q�E��1I��aV�o]�ϗ�z��UF���j�K��� O��c�a���JJ`I��H�{M�7�Tyuu�iii��i�}n�3ک���EO�F����u�m>�����>p!I���TX(0&;֜�)q�Q����e�"�U�ڣ�o@��-�Ri�>$�7��W�bA���"��w{�hc��
�z��N�I%��c;�	
7����@>g,2'J�dYȩ�r��qss��7n�o���y�Y�ws4��z�$��������u'A'�U����8eJ�k/�A�{���RM6t��2
7u>?����2:z/??���t����+�Ю<��,��b:f��^ʻd'�GT����s�Vx��	��d��<.�5V��;d��҇]��b'{pu++�Y��ގ��xi�2��H2.>�~�Q[��\���>�\��e���<��wX��?v2���u	��8��r/�.z{���'S�y%ڹ�9�<,_�(��R��̽��O��'t�;7�,�]�F�[���d�e������Qy@j�lpE�wQ*��.�����HQ�3j�7Cz�H޻̘��;&�c�g`-Tt�g~}��%|Š]���4p���J-�T= ���016�L\\<8���m<���v�r�zE4:/Qf2�����>�>��*0��RE�,^u���B�4�xo�6)|ܷ����v����O3E$�Ґ���x_2΋ۀ�ibY��jĴ�τe���m�P���m���=�ٳ i���ru��M%U!#�����8�?w�9��J��P�FQ|h!�>W�P1�-*lC�I�g(��I���&t�7�D�R��u�!V���/Ӏ6�lO�W��{^�k��-4��'r�!ݶ�����m��|��׌����X리#�_B�=k�%�e�z���~<^B�
�w`���:���ee �)�Y�{�u�{-��'��/�{���'>yQ�l�+v�>��6�e1��'3H���7�o
:�?���t��LO����I��D�������K�V	�Ǡ{C4tL�wJ,�tK[A_��-�ｒe�g>o�sX8c
��9��!:R؞�~f�#����R���vm���3���@.���9;F��hۼ����_�~Rh�C��)Y.%k��%���\y�].�hU��N�~���*-�r�4٩^�]u-�
���`���������x���W�8��nG���xB�0��e��z�Fj�*���������S@8+ܥa˧����������2�o���,�������-\]��.d�� _�L|r�;BU��~}%G�tE-���5@���@��҇�TV&�������-�MU	������_���9�z�y��
s����UN�y��OTY��GY�I��qFaJ#��$w���Za��o4O-#�=#�|�H��Ts;�bVªwp;��d��rP
,�9��:�l��B��������t���E�]^�d!L�?�w�LL�cH����O������u*L:T�>k��3�Z.��:]�EV��7���c��
��!��F2��Ǩ�=ݗ�-|K3d<�g�[Q���'������a�_�_6�^?�Q�_����'��T°2�VBCC��U����#��=�6<���=���h9�\���\#��!�9���Ā��T�����l�+m�ڡֿ�i���/@��GK�R�C�`�g.����
�r;��$ޜ��a��PPTd5)�>8��z�F`�|�^�/x�.sywK<61�|����ĉ7���y�|����#Z� ��=��&���mG����̺EU2s������yM���D�#�Kn���>o�P"T܆z�)�/"Ra0�'!��x��^�=ü�	(dt�gދ���$gQyxE`xx�낷�?�::�/-]a���ҜXu�����Љ_ >�Lz�1�5&�KP�m��u��^Մ��g现n��BJ���C��0u��:{�3e�(�uV��g65�s/����;�]� >�Х%SEEEk[ۼ�
����D_27fJ���)���KI�(h��$a�g~����7܎��r��UW?��@Ӛc�V/dS0�hZ���!HF��X�η\J�����[�m�KZa���΍���(i��+Q�9�88^���4�W�����y�(t�m2�����O��;�W����J��������N��ͮ~���������\>��(w���?���(v�/��۟i�RWL"�)"sʃ�r��������R�6n���;�=igz.�;#b\P�� eh��?=M{��ܿ�Lm/�է���]����L��?��	�3��P�ZZ�����.{u�3}�<_[6��z1$�78
��E��!�J�t��ڛ�e(��j_��UZ���l��VO�0��V/#�/`P�s0꧃�5�K-������T�ia��\m�
����V4�'4��xq4�Ȥ^�>=�LV��֊�W��&4zbC����<d/���t���>�_��T��G)���i�_���w��J��B�M%5�S_Ҥh'��l/�Tu�:x|o�eⅾT����g����1r�
i^��}$J���J��	�2U�[#�Q2]�	滃�| �u1�M��m��W0uqEe����b*=%V���6�D��{��YQ�!�U���z���?U�3u,/�Ol�=5����ac}3�GAS��q��V���A�#XC��ͣ"��3���!��VC;S�'�O�����z��aK�D��3rH}Q�I�;��{g� �G5'�`͛lEM�-���J�����+�+(D=�������.~岇�/��g��AV뙖F���^fCw�,(�>��-߉=��Vk��T�A⭭ˆ�:.�u��0�sˣ��ĬZ�'����R"�H�^�j���h�kr��dc2p|S��*�����~�el'��1ۅ��V>�]�t=�g�"\D]hP���F���>lR~���#7��u��>I�����[�b����9	�Ѝf����Or]@#� =�u�C�C[���"R]�D������b%�!м��p>��	e�G���Z��	�`��t�����D��V6�p��H`���W����vC�@�Ao%%�l���T�9�*�9�5��^$>�֩KP���4��Y�F�?�_�)6�5Y�O��J�����Y��k^�i� %!�,k��wL�Ԝ��]_���y[�7q#y�����>���\h�=�q~H  Ӷ	�Q�_��#��(�غxc�?|+�r�@x�W�/~{�>}� qfilQy���ә*@�	6�a�m4�)��HO�����'[Y��\�1���Z�W:�����av���)g��d��Y���H!�IR��C<3h�"�_��'!�����<,TZp���p�W�X饊m�>�y&�x!���ˣR���i>����R�}�z�FTU9�$?A��I�����4�3�qs�䐮6f>*/�.Ћ�hGy�ۚ+��c0T�}��8*Q�u^��)�s�ߑMM~��0 +��sP��"ߴp�&_J]�_�X��>gg'�$��^\\��e�Ɨ���w��s��V+j�{�"��!���HBF�~ۋC$m������b`�r��QKY�Ī��n�)��}�y'{F^�{�����&0q��p&
w[����'�m����/�q�\.����?iĸG�#�{�R��o�����!~rF{��XW����&a��'��w��$̟��S�A�>̈M��j�T�,Z�q0.��ϧ����q����T\HZ�Ԁv~�W�j��OMK�SQA
rIII�F|���.V�-V��$�%�h��AB.�`.��q�Gۙ*נK���(d�p���`%�e��&>�~D��aLF&$̵1T�(��J���������=��	+�4��~MiQ-GTQ��=�_.@xK��h�����/t$G&7mZ5�[�k�l����ޝ��a���y�^�?�֚Z���t)�����_�.־�1S�i�A�Z��ׄՔ��k*�5j�\j�ڒ���ˣ���%�����Ѐ���G��! K�����[�G���>�����z��b,~K�y�Vk*�h�Q��()�y�J:�]�M���|S�e/�#��6����"-nմ�����g��������N�6�����|hc�;&����o8�P32�2{��6x����W�����{��:�[�.��=�ɭ q�P�~w�x�����Of�yj`=r���{v䃂�gD?�l��5���554�3�8���y���I)���L,����ى��:y����:p_>�joW�'�IF:ڥ�1$����I 1$m�]���W��T�$��PjA���Ҽ���^;/�%n�Ҽ\[�u9-RwX\.��-�[�������=$��`u柅a���br@�day�Z�\)�����bIF���R�w�.B������d��&s{}@*|C��i�i�}m`��ߛ0׳�:���:��U%%����\F��Sked|V7�>!|#~6Kg?�P鶡;�'��2�W�8?���\���oATF���k���'�{gEX �w$g�Iz)�6��oM�}���P���t\�m?>L}��ɺT���h�ݬ�m_��	E����4`�OCr(�x������m��X��_�PgJ���̱pO,٨_:Y���'h#R`�I��t/��N��,�6�G!�IsU�l9�U����S=_�w����}��.��[Y�)@�aL	 ⸵ۋ����=�\�=к�7�cڴ?��s�ۦb�B)T�U��^E�;���ǲ]�ML�l��m1�Hv�d���Q�A��s�s9>�҅�K-U���X�>��νCbF<��D��x0�<}��t�d�e])�)��.
����a>�hJ�"+ Z��ɩ�^� h�n0�j�&�g<A��-'"�J9iƞ���a�J�l���Uq;��O[�a+ГT����{dB9����ֵ�d��B�	�K���+�ꕧܫwvI'd����Zᣉ����}��r�.��O�:h��P�n_�]"}�}.��a��b��]�A{誋�B�o*EI����C��Ba�9���ϳ��|3���6#���j	
ս5�Q��:��ǫ��8��^v���9�1�G�ɏ���6J�\HM�?��_	�to��] ݭ7�6�j�&6U�߮'P����m~ȝT+�U�HY%nnw�̵Iû
L+�R�[��zxp;�[����w�W�
�ĸ�I�14���v{���L��f�VU��e�W���}��t|��ܩ��ˢ�ƯR�~��Z�*���/���~q�;؀;b�M��a���a�Jw�"os�üE���I�$#����ҝ|,Ml��KxCv�H��������.��2���-�-
h�dUu{~������ʵK���U9]����ǂA甡m��9�=׋�=c��T���$l=�Е�8^��+����9��Ꚑ���m�>�k�(�(��ݠȫ�쾯Ƭ;��Mͱ}�õ_�$J�M�N��K6`����@#�є����є���f���L$eȸ�����>*�۹q&«贖���x}�
V� ���������M�d�dí��{T�V���DK_�8HB�Ov�rjG ʻhlX�a򍕸uC�>�fY��G�n��h���:����^��K���+o���l{)����Io���̝�����2:9�`&'7�rx&���0�^\;%���_`c�c{��̇�dZ������$%��sWq/��iR危���ى!�z P? 6���F��j���*C�H�?,vC��GLw���K� �埨����9y��a�j:4��s��Yi��d#=�� t���黫Ɵ�1�(�f$�<�X�<&����i�qm}>@��L�rM�B���*¶N��� 
��^�ęF�|���:�؅]J/���!����z6D�_*K��8�렞w-������<�CNǊ���^���ۜߜ��=(7�=���W�S����nuy1���n��� O��*I�".���j�!O6X��.�[�9ȥ�c�A���6))�vӧO�6�h{Q���'��V
й��}��&��Ѡ��%�#��A+��TtttӵV䤤�)�5P-`��<;U^ee�G/8�a(�ؘ���,?3V�����;���VJ=�B�'���Η8�����Tј	�Y)"˯�+�����޽Oyj��q�����[�+�1�c�����fzkvOA��<���!0���Ax��t��B��kZ:�r�%��F�x����QY	)*��_U��,��&��ڢڵ}@I�\���2A��ÓcwJ��V�ԃh>>��	����������g�(ݤ�xuS������K�U����"u��\Ǖ�3����#�������jNS[[�Z��Ů����l����Ҿ�;E���n�����%���10�s�q��b#�M�rwH_Oocs�=<=�}T����z@��z�v�xK���CP��������*ĳ�4)V0��jRgj¶o� 	'X�7��<9���z?1�$�&�5"JJ���{Z0L�C���ŜZ�2YG$rU�w�^��Þ�m��7?
��=�_�J����o
�+0R�K2��om��8�;���}�K/�*��Y�#�j����Z.�C�h�[��&�m��*����0)�
ein@� ��+�d�1����j�h{�P���#��#6��P��x�:�s
�f�u'?�����8�����zŖл�����۲�:-��?$���\�3i'Z����SY�p��P~{�x3}�n1���y荢�<�O=�v���A���U�U�z�O�}�����&bxwiY��e�@F�kkw(�p�i��|���D����P���}0������.x;�В�Y��5�ժڒ��#���w�F��4��b�B���cCa �i>�*~�%�a��U*�ܖ���jGO,����C�D�q�虿tZzzIII��0��OM�#��}�NE���!z��d�r0�N��K�0=��� ��FO�7�bTI��L+��ͬ�?��/d!�\M1 ���2�JғS��~GI�^�����rƣ�"�濈�X����io|��eaz�(b0P:U��`Y�q����~�!�W'E�V4��%�z��7
�)(ۡҮE�W�م/u�����.��%��/��0x���op*9%RvB|'���r�9嶈�4�4j#�4���w�ՠh� �>�*���|����a����[Z��׏��/خ��PSg��Q[�u09�}yW�r�\�u�0����=@>߮��iN����Fl��}_A�L�Y�U�Ԃ�J�S��E�T�p\2��ȧ��u���7���Z�}�&~�j���qa�~eh�����m"������@�8P�Cmmm��fꪪcp�:����eJ�q$.�v\ɝH��#k�{ېg��=s���U+����)΁�%��<dd\oљ����8�-�Ӌ�k�k�R�$�s�O���
�^�n~g�ރ�V�u\&�v�_g��8U�f|1�h�YgM7�/���
r^�۸�u�x��d�A@`D~e�c �=�� �|o2ג�O!�S�V�X�q��n��q2'�Qy96t�XF}aR��D_ �
�����+��9�-����8���z5�O�/�8�� �k�1n��Ӑ�J���3� N26��Sj�"<g)"�nkRwfj����1�\_����BPD��,"��f|�Hex��=�����E8�?�G���Ў�c|&q�#v2��B|��W�J.;�3f�]PM
/��1�LQ��O��o�;\
��21.�ŭ��?y)H�6���$��F�ҵ ������m-�MȪ�)�e777��������Z��pcH�Zf�We�w�@ ˷׭���?�I#J.�s��A�'4)�ppo�e��M�?d�<:���;�D��w�S��E$0,���b�UUO)*�=����� �|A��Ҥr<WB������H��&I���@Bz�x;����mYqÂo���� %H}�>�{�M>��7�(�{g�޴�/z{��Ɩ���~�F`d�spv�SV;���h��6�)�!�U���鐍	�#H&33���w���rr����[�5
�������)���+hJ+�G��R3��m��5�q�+�\��Oi�S:۬�z>Tn\�U���*��#��JK���-�����k�U��6#����=6��J�E�
��S�..,]99���ޛ��}����>�������ςA�x; U��wo�ʌLܯA��P���HKO�n�RE̐��m��M�4�AL~�
���ZEj�^آ{�&���:3|6�x:��?��f��pu�og�%j'�K��j��~�Z/KҠ��M����&���^ZZZ����g�Յ�JV��W�c�;bvV�vjꏲ�P�o�y.����=�q����j�[cJ� =?���6P�M*I��մY��Ķ�3�պ��p��8��r;\}��b����)]̷7l"����up�[`�����&�9�>_eb5���Z��",�P�������c��Q6\W<�@��73,���揨>3��Nś�D�AD{��wJP\޶xT��rod�/��Z�t�)-{Twyf�΅t�����R�pߛ��X��Pք�wbKr�T4�6��	�ƌ8D#��.X���{�!�-3ӝ�H)��.&���flRùk~�ۆ�vK�����T�
�3w��~�2$�]�r,�&�6���qnUU�*�tv��~�~ųP}��M
F�+��6?�[�vCc�O��9� �.y�#��i�?���x	s�V	��`����h����\_����jv/�*�2�F'����!6�?3agz�x~�Xgsi�Z��8cl�����^̍ pl����\��6ۙpl���R���_�)�PJJ��5�$��\��K�շ*R���#|��h��u0���LG����>��ϩ�����ԠF�T�N��g��F�.�,�y�6��3���뭪?��:�i�3?�5i`�۩]U[���ѷ�ٵ�s�/��Y���	(����g����=d`�a�N�e�C]ȤW�9����V��8|zO��hs<;����Ң����*�S����9�T�bWD1�d|aA������8�P �7�v}y��}��m#Uի��0.X7�OK]�.Ǵ ��S����۾�ֿD����<�2���+J�eN������ǿ�oL���|�QW��C��fa|��e��;F"��G��%�r�K��tԟf�,:�^S�+-���Q��+��f�o
6D!oV���m-��E+��49�`u����  ���A�Lq���3M����k�;�q���2����Fy10Pĥ�OmM�c���u*�E�l�F<�o,j2+-]ъ�F'ۚ��LQ�x714���Wv^���\v@6ǽ�z< ����*��K4v�[�]i!�}
��c�C=���fuVN�OqP� �J���#JNd�fbr�<�7�jOP��,	����pWey����� {��mRH��Hw@T��o�I�V6v�KKd�ZI@���2^U�	]�����]��k!�騕]5̬�U�iw侹S�ٺ2�_�q9EB�6~�����7��kZ9_T���ɇe�,�T(x	��p��r����:@�	�+v����*���w/-l�JUm�s{"�S����=l�Nv�0<7�Q�� $�Zj�G�R�՛�a��j%"rrr���ZA�Q^[[�ƫX��<���)��񖔖ٻ����30b�/!���&�f6���y<����]����Dx8G''#N�
���� ��ܢ�X�3 Q�~����~����# ;�4g[�$�r�qG�S&#�p���˨���3Ħ�Z�$����BE�������`�/� ��>60��Xx_ߧ���l7ދhP�*�t���B���h�Ⱦ�v�d �C�����!�I�͜��b0Юџ$g�An��Ff'��i�N��̟��SS���օ�{�]觡e�Jy�;�J��+Mf[�^A2d���F8Oe�u.|R�yS}�gGm��%�V�'�c�v����p�:>upp��ұ�q~c����H!��U���6-��&��o~Ӛ�YeOO�{s��KK����أ>�
OL��Vp,�5v�pt
�3�.���ZvR�G�@��΁����-���nR~+I�.�4�݈�9j��C�Vۺ��n&��rK
���躗
�@:OT!֎Y6ϧ�f��5���wW�4� �S&���#�c�Z�Y�`�b���	r��!=��)Qr��l0F>�9�1��*`GΩ
� Ĝ/Eo���L7���z��e٣(�����lX���:�f� ��ݰ�M0�W� ���y+�u��O���Um�.J�����i;�ꁾ�	������o�X�ݤ�U��\t����z���	���u+��---��6@���J�Fm�o�e�&1��Sf��Xz]��\Ab����Xp ��T�n���t���x(���?�
��~/�02�F���Rg��6i�=�깍�D�UTR�wH��TQS)?;���p?>�a'�B�'Sr�(�楠]0Ƅ��VlRy��3��2�߹�2�k�#~r��,Ƀ�A7���b��Ee)'#���0N�KL̰�T��o!~	��3���y6gm���hc�1�V��^�K���3��lߨtr��������&���q��\�k^�1d�d)q>��}( �M�/sJ������Qo�29�WPg�x��l��K�ˬqn0���b��V3��BR�Z+*Q�fff
Ò��0���;��0m�w�7���	$...�u��l��g�����˕��� �[�p�S��. ����\nz�Hp��͒9�� ��%�?AWU7=��47��3y'-�%0�`׌���1�.g�gD��kCݤfaЭ�P��w��/�[��P<�]��>�ȏ(*������vZ�H�{),����ͷ�B,�SfD�G����
��4D踠��<Gds�YŒG���hz�E�+��2����C�Z��?:��Oe�^c���H��Z���6�].!�D�[˭�De&2�s54NV��o�I���_�ְ$��-W�᫑Ƶ���t��`s|�YDY:Y_����@hAuI���#�hw�Q��>�UU��_�-�/�!S���|���l	_.y��E��x��`�:/v�q��a�H\Ê�"�"����zVhi);k��п������Ϡ�{q��h4��=��X�h�G]����&ׁ�W@�l�=�����o+�q�_��|-s����(No��^+�K,}H�U�qF�!4�ot���M*�Gh�J��UZ�~G�J�e�\8|�d6�X8F��������f��(ڇo#�{Y�
��� �jA(����z�Pw�fOtX������u�n�;K��7�Y���;v����	���T�]"����)Y�P�Lb�9����g?ʜJ�>��|�3�����t���⮮5N��s�*���s�/���X�G�3�8y�)m����Zn'aؒ�үA!���z��=��y��Q�Q�)g��:?1��{��W��x-���nΆ4��fT^/)1��Rn�GE��Ï�[���{�հU<2�~�/;�,qDr��z'z0��EG�������t��lB�O/�ᨙ�A���U4�F:Ih2|��%ץ{�����@�<�����	?��z�q/�d�2qY�	nyL��p���/��>��j��+]�ů�M�O�g�Wƒ�>}���(s�;��:����4\H���G�'�bN�n��/��YwDv��N�#��'�_5��A�Sn��,JVUu�H܍2�y,��4��3�0�}��G3@&���[d�y��-=/׌]'P�gg��'Ә^N_�R��g}S+#g��
� �t;�y�Ob�A��>�l�����ߵ�^����P�fl�F�,���r�(w�h֍Kl�^����=��������
�;*ko���H=��+�my�7{�Wo\]����1݆]�s�f�@$�߁��K39Ƞ.{0���w�e$[�cj���qtt��)�J�RG������Bh�+�1�?u�4<r�嗳��K����ӏU�kk0�|tv�v���#;++�"/.#�Q�E�M�E��e�2,E �/�}�eS�ܹ{����&��ɪx�csu���R<m��������:�i--��	��.�H�U捘�UW���'{k\�ǁ�S�-�|0V��3捹 �~?9I���I;���PMAƘ�F�F�VXX���_
���T��ӪJ؉���ؖ����[�G�F�q7o3>ݽ�V 3<��+��+��~a�,��b�T �̟���b���N�,4��v�i�4ß�_P���a�����s="K�����BV@��C�o� ���+|�m�b��qÃ#Ƃ�`+���D뗠��|��P��+S�8 �l���F�U�zҁ5���Ǎ�o�D��.~A����=�Rj��\�[I�DG.��7�?ή~ʹ��(M �n�,��CalU`b�����:$C�*
�pv�.�����e��t)�'o�S$���pp�l���Ж�I3�?��� EJJ������#Ģe��R�x[R}���vx&Y������Awiv�Ul�@K� �@{`�D�_��狘n��HQ�t���{�-O����e������ J�����lTd��}�fE���L{�>嵃�G���y12����n�.l��?����+�`��l?	"B	��6c�_'YT�*-��ʵ^�{�Z6�t$/x��#�M�?7uƸYF�r22�M��"�u�r����6��3�~����LSN+w���F>�h/z�%���_t��
m��;uj#��ة�<�������Pay�z�,h�������U���.j��w�i���g׺�4�7�M��\�g��f��>�ޜ2���x�(B���{=v���T9���֔��/Kz�?�g��2���}Lf��O����ȎW{!_��0���btP��x��$dd8����c��%�n=�y�Q��\@ �򩚆�1Xb�5t����e��<}szff`�YiQ>�O}W3L�!�$/�%^XQ�`��G޵�[p!�����S��Ў����ՖÌ�ꊓ���g�݌H�����9rW�ē:�a��4��D#J�û♕�m���������i��VDcC>G����S�('k�#�������Jx�0a��I�1@�3X���@�}V�n��b�]bh0��S�m�Ӓ�A*��C��{->	�Y�kYI�-^�����(w���;����z!��ak!��� H{]һ2��\[���!/g$.�?5�kؽo*l>�֐!^s695�T��,��<	x)/(>�&��e����^7��پ���z�ݰ�v�+�xk�#���۲�pq����vS-�(㊷6��TV�3�*�NF���Y�gN��X���Q�{��G���!��R�Bw��.o� R�~�ʠ�?��	���|�������ky?�ǽ���Į�Xq�iU����|����Ia�Ba�������R�=B��R��}7en�VF����?4���DH�NG#��4����k7mF'�9�;6NN<���ϹMZ��[ZB�q~,�Q�리�6����`,�d�1K�m�J�,
�uXc��ѵ �8ξdQt�9l�%%���6F,FȨ��]�8t A��ƳWl���}j�*��M��V#r��GOճ�T�V�S�`?��mG�׊�K�$s���}X@[	�0D�p/6sǮ�N��,�HM!�9����Q}-�θ�HX��9��N��Y��\ؙ�=�"��o?�6�޳�[!5+ �HVN� �o���0e�Tss�O��ͤ)K��jj�||؝kϡ�0���JMaMJ�[<w��)��)gaS�^���M@�5���e�}�>��F����y�Lh�s�I�'�*����Y�����+e@P����ڑ�;J@�Ÿ͗���������@n����3G���ǋc�BĪ��z�m:F����K�53�����J?$[^L�k��8�T`��N����Jj���~#I��ST|�_��9_R���`Eff���N�MzK`�v3*�����)it4=/
\��O]ks�]qSԼ㖠.ݴj68������s��>4��G�q� �S���<Ԇ�y��������/���/�y9r�_�o���e9�/���M+ۃn��p:��iu*ރ7�b�E։z����!���
q�gy�[��+�f�Le���*p1�鹯�-E@%N���Q���3��4�x\�E2ҿ��%ն��A��i�NI�¹$�ĺ��CxM���fO�|�'��ؙ;��͍<�,�d�#�r��&q<*��?�D4�Z�H���}2�8RY袇�Y�c�ZW��Tb�A>}N�t���<��}Gn�1�zj�>��{m����hûF2%DL
�I��\m
σ��|����⨥�=.�����%;�,�A�ӟ9A�&E�(**�TT䶴�om�rpp[�5ī�m���y��s�P�hS�S�jx�yM������^N:�g�!s��ٟ��ڻ�v��ϔ��ϫ	� �^B-�A4\�}��>���/��?Z�;�pm��y�$Y~��یx�@ {��(��c�Gg�H�U�V�ȝƅ0�	�����g�rR0����q�ͫ(��c�)'�h��[�zc\�y�l������+��U��u��~';��y�k8G2��!�G��� 7�S�Ӟ�S'�NA�!QSĿ�z�\f�u��pkL5'���
'�;Ha��c���:���as^��v| �v��L��S��}���І���R���&��X��<~!��Mbcc����}�2��>�J���;(��?�n;�ax8��~~|�����"����{�e�"�sQ����6>�����Y�M:���ୣuL�R�գ�]�v���g ��@�&�"���Ӄ��B���[Gm��������BTR҉���3���?��rkbH����MIY�V���^�1G[%�P�!Rsj�]�I��h�.��x���ԅ��'R-���O��X�@k����j�yy����fq�����&�]:��`ܮ�m�A� .�ţ`��q�2R��2��A�{�����~�H��5�d�C1^�+�GR�ӵ�Z ��a�#"J�KW�K�� gb{�ǞF�7Z�Gr��cKp>�y_XT����Sfu���\�g�*��#*��I��|ƶ���ԅ����ޙ��Ļ�},�l�ZD)�=���쩐�m�r;�.bSD��g�cl��LLŻ0�iJ�%�:t@�+���K���@.+��,P��\D�4S��O��<�y��6����fV�����ے� ��;}�s6��7	�/�찎n��|�4A�|W�A h��|

��+�ηw��C�"�I�4���T����q��Yj��t y�|_�tB���UZJ����(trrX9wco1�*��~��v�34TNE]��z��,?�fͪ.&�*V�©�Cֺ{�t�%�,��q*��m	�m }xx��ݝ�T���N���(�h5�Ǌ�������q�ss���VW�M&����c�R%M�:C����6)���³�A�E�R���2e4^rgw�<p|)DG��������ɮ���d#��|��eԙ�I}دH�:�N{{�Ʉ��o��)���=�Z�l��::&�a_l^r&S22z�+�y�S-�+ro;�J�k6P���X0:�'�x��7}���9��4"�SHU�)H�8���(��rP0p��W����N�G!A��a'nm'6iT*0��`�^��7͙�� � ��C���`k{��09>^���\��D��kXPp��}�!��\/��m|�
i��~�qb�c� Y����i����A��l���L�
U��B�g1�\D��ql�>퍚��m4�v5�[���Y�E�ݝ����$��4e�\:S���ˋ��c���p����֦V��v�M��֬;����	EQ�(�ڵ���=R{��A��������]o�+�T<�q�}��9�t��Ӛ���<�h��<-{�ک��������UbЫf���Mb�R�%^_�z$��;t+n�l��YP�0�h^�;�Lī�qST��ð �I���;�j�=Z���F]α�7ԣGarF]�&9���bw��}TIH2����Æ���SR-�3ʌFߢS�u�8�j�aE�C]�~�Y�ʟF���R��y�0�>m�{���Q�a����]�0�'�\�u��n%4�o�JYLAb����;>�������O<Wv��o34:
��&�1C`ˉ��Ż��d�<��n���A���Gr�'��w������(i�Z�#������
8�s/��<Ή������%���=�*+�hc���p���
���삂0,���/M�*�/o��=(�z��YY�	S	��ٰq1�(�-}o@��o�r�߉�,����]�Z9�K<$Ϫ�K}��BA���2�%����rY���ҷ	k�03�R�,��R|SU6~�l���r��_�_����.����}���uR���	��^���q��*hd�������:�uv�����~�9�;�,?���xaa�V���ٿ���y\�ф%7׌5����C�{��z��)��//}�}��%�>�l\Oy��1�э���%�ΌX?�����
,����p��t��o�.&�:(���'8�^TY4�-Q��X�N�F������[����Ҏ���!�_ip��t�<��_R	g�N�)J¥ִ9=�`�V9�����9��VΎ6�tKX�76t�7ꢢ�'&$�mP���}���M�㌜��[*�lq�NfswZ�J���Z��i�A\�2D��+Vfd�=��|��kӾ�1�g�Й���<y}fb2S*{���z�1�b��78�=���H�0[��r���R�IG�,�u*2W�Z�rM��:@vՖ����Ӥ/�0(W�^T~�"n$�ހpbz	����u�>�[����]1L�CBӿ�صhʲt��%?X�XK����X�aj.�T�����ރϘ��ƽ�\�:ڜvz�dK�xmb��>!�]I�f��%'����a�</v���(k�ХSY�W�D$$G��7��uuiKJJF��Rq��*0�`���R0�>��߈���=v��Х��)��/��%qB)�����y�X	����?�)��lM+�$r��1�(�&?�S���s�P��a9�+#�'�`�R��၀�Xs�t��J6���e��&�E��[����Veku1Ph!4bf�S��_.��'k�M1+��w�@�S5��C�o��l���?��}�JiK�e{b�_�H^x����֮P���Y���r�t:/i[�P�#ݥ�ɠPS}���j} �N���n����]j�S����mʟF��4z%-���"�97�n���q�eT%��r����%W��ǌunᓓ9��U������}�L+/���\�7�	�*E%tت���{�ӏN��ξd��Md������"��kl`U�I�L4LXNI@ƘUP�<77G-bX�8qa��y{4G�u��<�����;~��.B��&Z��-o$2��V` �.�0��u���񖩏=�J�g����o7p5?�9�3CQ1��T�U��܇e� |*|�J�ቈl�zK�K1i/\
�ۨ� �-6��h����>���"��%s�r��>6����~7����?��aD�g��7���ZZZ7*;3CV\sV��Y��1	��V6�!��ֵd�>d+uj�9��Wn�r�,����S�M�*��h�?���Xsm.�@e�m�E��������_������8H����ҝA]�6��t����Xy��Nڮ�T�edd,J�W���F�
�`@�K�+�D��]���h--��Ig�u�̏�IʬR<�Ʈw����K�ﮤ�[�����?��"�֠W�r�af��!���Ze IP3�t�~���6� � CCCo,3�NC�[���<�Z/~�X�͢$����7+�����K	��"��e^��L�R�{�_��?�|�d�@�����̐p��̨S��[�ިGqUb�K҉j�ާ\X��~���
Q�:}�.7����U0���̗�$��>����J�ܳ\@$� ˟fŀkL��Ŋ����M�ggw���c�������`N���=~J��W�1���}2[�eN-�� =S/��%��e���g��[ø����\"��kX�\���C��K�c���0�K�:�>^^m]���*�:Xd'�Ol��$;���^��K�eZ��#�z��Q��-�Z���#C��V����9�W�axB�w7fkV��*�.<Ӎ\�ո�� �x#��$$8z��Q����j������
�*�<(�M��Z�1[ �\�FD :v��y5J�b�4�x:��߽(���Sf\Z`ˡ�Ն��(���D�s�j��d�(�?U_�\�|�vN���e�ʁ�'z��UP��n�({����0 R��N@���@g�Ŀ��G\�/���R���L�k��U�}��Kn핱�S�FG����}�~�r�Ô=������%xv/350S��LW{���$e��y�x5>���3tGy6̏-]&����b���ɡb)P�v�����W	+���%VFZ*~�.�w�q⍌ �|�~�'���fX�*Ky}�$����ٕ�	Ҝn�����>�I��Bsf�LB�5{����^ ��B�Z������/����-�&:f�O*��F|�����n���?H�f|�6��l��W�rCm��=�0al�<�ۿ�jO�k�(}�r%�������ŋܲ�t����ϛϟ#!!�  PX[��.�v_p>}o���YOB��gL��J��Қ�G��Ѻ�+t��܌&��)��$�Q�(}����m��]����Ja���g�S[��<J�j���"k��32SVL������Ɵ�Sz�?fi)�N��}���P���k/ �q�p��O�&�(�3�G���|#�=����"����j��L]�Ɔ��%w]��g��{���e|f�������߲p/p�����P���O�}��_�B�V�^U�M����{=�����S=jh���i�UUU�{�Z��Q^�M��Wf�z[ 
	�mP�#;ܙn��vs��9�6kf����Fqkz&��'��\.���hc��ґ�ڥݶ�;eC]�l��2�ؗ���� ��̽�� ���S�T+��2Vd`�,���eIW��0�%�`(_� F/���칳�^�hΜ�s:�K�޾����L2������c���q-�{[�/q��&Ż�6����5=���o����;X�y�}�>�2Zq�ԏ�k.�Jy/��5!!�o���wuݽ���8!�H��z<%�+"�ڤ���f�����I�w���Z�����ę�{��x{:���7;-C��Y�N��+�g�H���������[B]�`��������N��2�X n����-gm��_F�Թ�|q�Y��K�V�לj�Z�Ã1ϐB(��#2�t`'���7�ς�VS���Yy��{:.Uufі�j�9�;��fDr7�w��p�SYe��չ[vj��s��̘�~&Vm�m"��8��O����̀�Ɖn�__������)���_x؝~��q9�4��c�L[R.W�{p	^�?�5P6�*6-^����&����qm�^s[[��*������$���
Yu�܂2mCv�����n��^+x�����N�e�;�U�19cܬ�g�bE�����?M�x&"S98��w�,.U~�s�R���?�V��i��"-�s������ J0{�U��9jGx����{y����x��A>C���0��VE�I�p�#v�C
�G��<�>n�7�`G��H5r�-�i��<mcj��H�Y�����+}O�^�/ŷ��8j=�;|I/jn�5l�;���|Ul���|��*�K�7�a��Y�z�Ɖ]M�F1a�}���Q����^	~~��$�k��֝�����-���ȬH
ޖd��f�Á�)��Ǘ�������{4&�����6�\�{d�*��͈�u�� Æ��cx0|��{E~��R'�W��%�xĻ�����VX���2Ϭ�����\\��$��d@F��w�D�e�<D�>�b����]��E#� �T� �㹮�΂�a���[B�����A�҉�� [��:�ˡ���@{;��������\�Nݝ���G��&&}���[`��[u�Ě{�d�{�dX�G�-.|~~}d"tխnz|T����R
�(}����U�t	����@vN�ć����ar*��8�Y��B����P�W�;p�3xܸ����'CBa�a���z�xBBM~8}���ӇYC�U���ѹ�Ŧ�qp��yЗ�a�ttu>���
\n6?�}x	�%b�^ˌ`N�(0݌���A7
C�Nv��gꐈC"��2��+QY�{��HM+�`_�?�pI�9�6���_��%s)|u���q&w%}���뢉�x���[�jk�ji�^��RLp�W��xKEK��H�"!�B�����Y6��}������32�:�U�>�-������l'y&��"��3Ǣ�z�6o�ҖҧZ�7�<���5ʚ��f�d%l..�����t��䑊ݐl���IWǢ��ۻ=(��T5�o�?-VmY���(��N�-Ⱦ�@R7׆Ob�v�ş��M�E,�	Cu�ה���UZ�s�V�nK�{�v�O{#��z�c�Ľ�	�H�3���E��}��VI�Wɲc�F;���X2�绻������6�����<�h�������*3،�ݻ�[u�&dP��3�Ͳ��;}�MO^	���H����@�6ʦ�����y��Z<@�q�هWE�f
Od����x�b�92~�~�{��������H���N_�^*�"�&���٫3��_c��r.�OnX���=]F�!���!͖^fه��8:�꽱�r<7^���-�$�U{�z��$Ht	���T�����j.2cF�X�$�����=�ȱ��f����P8���l�K��ￚ�V��	���)�fz�N%PBfj�j�{)>�^�4ϟ����D���!M��>2Q�PG_�flD{9�شn[���xxV+��8#1��"T/dI���j͖�J�cRn O�ئ�A�6.���神�k6O�W8���k���ՙ��~��Ƈ�j����B�Z|/�7�Rw�����+��`��ȭN�hLEˡ@d��O� ��bc�O+6Þ��ppZ�{a��vS�	t0��.���M���H�jKN���9�e�钦
���t#�On~_�L)c�a3,�Ԃk�*�&A��|rɡ
��Y�W���:��Ż��o*��`�r���&����� ��v��K���kk��S<kk�b����2N_I�� M����~��i��5 �[�h�;6S�\2����-�w�P��#{��G�b�3Yj~6������\ �r� �c�s..��Ӥ ���גⴗ�o��V�-YnPdmп����MM��Z�.�8',�~o�YUV�M��E�4�Z4$`���^�^��FȼҀ�V�
�зP�lݭG�i��2��KwC��w��a�4�M�2�܇e��\R�2z�XeA�!1��Q9n��;eZX�e�2<�ߴ�+��S��0e��,[����R5;s���b�?)�F v:W�����4Iqݖ)_�fa:HZ�T��_&�x��ئnLˌW�*(Ȕ����%�U�#LW	)����N)'����?V�KJ�S��$�VdءT�ie�� �Z�Z���o�}8-{��~N�hO`�
��G�1%x�}x[CKatl�7�g�(�5]�Ѳ��Qޕ)S/kƍ1KP��C�_MT�!{̬
���q�m���y&-+�+!�<G�{�
�<��@O��#���=Wؾ���쩳8�8�!(�� �r�d�����d˿�p�p�����,7��.��ϰ�uzyry�xjJ~;�τ�2|��u%�dQ?f�)�43n𙛪�NӴ��6�؊�[i6��Z$M�PŽ3��'	���?XfNvV�A4�73�~'~�n�Ln/+��_��eY�]�)Oo�3��jnQY`~ǝ����B���K��^8��U�)���z�����M��sd~8ډ�r1
��㚿DE5Ϗ�K�Eĸ{{�Ubx$ҧ�ٞ�h*,���]618��	En44f���ؔ�J�ݞ��	�FZ��S�_2���N ����'Of�U�I� �	mc����x���w��|�c�+О��>��!�k�:�r�MFIqO���Y�9��N u��s�\s�����j�/8��_Q��ں�>_��>���47IUqFSDFL|�E���7]����mA�%�~�H�zO��l�?2ftw��݅��gN�~-j2����	���-,ذ�V\�kv�a�Q���ǚ�����Q��|τ^������m鳶��]�	 �x,���=�̯���C���)v[�)�t��Peݱ�����7(����W�˂�[��-Mk���/ �*�C,����n�6�S�tM��B�x3	�ﭚ�v�h,�m�=?ޚ�I�3����$�R�J���f4�TT��U�W����=+|1Y�5i�ҵ~~��5.R�R���˓y��"�z�N���s����z�eLa0_����Ymlt��k�#_^cI�Ew�]� uK��پ#�+z1���l�.�Z���1L�܋�ޣ<�ssN_cbHCCCW���ST4)��w�ɜ���	P3z9_�)�D�z)�����E�#����>��\YY� ����-=�5A�A�����VZ���a=��f��t�McO�[! �Rdd��kf"��/�v`u��Ua�ၷ����Fs�b�=��M_�V�[=;��!^��������<y�=��ȧ����5~srB��O�=��r:F�w^�U܋9�{>{^�50î�>�퓑�D^6�\N��Dκ�pߴ��������P�v:��v`�SSxԈ
|F��n=�fڻ��4	K5༫�~%�.۳�s%�ū*��H�yQv��T���KU�gg65���Iݜ�+�� ܝ��l��-U�7�C�m�D��V�w!�b����a�ryY�v9:�<�C��FKpr�oZ6>E��Y��؈/�I��{�h�v�6Wl�ׯͬ���8�~�2�'#;: �U-*��e��ޯ�Gϋa���iqqu��^[�l���Z�G�����(C�а�۸�����)�+^V��a�|���Y�{M{�^���j�z��G���������>�2o�����=A�bN[�"w�g�k�4�����3�	�	�cy�����:k����5��M-%M��J��c0C��W�t��0B|�xN����}���M{@�P�����][�RW'ٟ)��+Ӌ:�a�kg�g@�^��Wk���˺Hm���[KbM|`",���X��g�ݸs2�8
��Hy�C�Z΃�$�|�F��ed��;�*��B����?uMt���"����G,CW������>����{v*��ۿ5�F� �x㜾��N���J�����~�.���N/��Fu��b���5�NfT{�[cU�M�s7��z͌�!��M��2<���c�N�܄V���f9O���%�ox��xd�<�^��J�^�I)����(�L��2{j��ve��,�VN����ڋ����m�j�&�5�b�R�}�]�ca0�~1'�bՕ96�ɫ�����b�=/醹������{4�N�A��(�z6F���+Ŕ�ػ,�d�H>�1��m��伽�
���ـ����.���X��@��kk� ��794K&��2;�X� 0�U�E���fWvAkk�ͳ��+�F9�%!�Y[����
t��~�B�;l�����R�&N7+���pjN��V29|���W9a�@��tu��`����4<�x%� S����U|�X���` Q�DU�B�5O99ɏ鞒����������t5Ȓ�o�SM1�璨6�<e����kt�m%�|�i\Jаvt�B�@ҽ� �q��7��\!T"�-�̏���s�_u�O���d?uV�Q��)�鲖� ����<7Y&�0eF�rqsO��EΌ��011	��8��[`��)�a��i"G7��M�
�J��oEH�Ŗ>Sӳ����e.�x+���64;�גFƱ���:<:�'�{�q}} �e�ٞB_K�oՙ���;H��_M~�	�l�I�Ž�U��l��i��e3Krl�B,��2�U7寊�Z����͞����f��t Ǣf�oA	k����3M2֓�ojIO#�_���;r��0�?�$SՎ,}Bbz��X�L���g*"ݷ�1t��g�~,
����y�Q����(�c�/�>�ri�O�A�Br�u���e��IJ�㦚He�����T$Ǘ�r7����ݔX��˲�YK���9�)�>��KM�O��7�F�[^����f\�$�!��nԹ<��ɞ�(��nQY����������D7F���5pz�o��w����Q�&v"�GǑ��혞�]�7K|H�<:Ypc�R�Z���T'w���O6��?�4ۻS�o2�-R^d��c�%�꣱���%��9�^;���0�~D�����d����
hq��������V4�uA%3漉ҙ�u�|��eK��m�'5y� ���*�9d�Sn��h�Q�RZ~E&��1QQ���{~�,9N�#��n~o��RZ}� �Ұ`���dTga�h�Wb�=��������*0��k����x�ن&���}�4UA�sz�	dq~��\�vsd�{[��@䎴f�>��o%1��/�\>���π\��J5�p�4Qg�O$&ߜ���`��]&�5�7

xX��32�}�a��O�jل=c�t�_��� ���J�W~�3O�	1�y����6S�9Ho�82�������B!id,S�?�8"�K�!��}�T���^��L�9�K���ELB32���FK��p�8#�T�O��GD=M����X�پP��XmJ�� WۨF��9�5`I��'�����&�{A���'���vM�qCW�2Id��͑P\%����2Y9��98_с��b1W~~��o�a
'ͮ�9�¹�h��Zqs����Z��Y�̝eo����ʝ����x�>{f)���4�0���x�Y���M���+-B	���w4�S�C�[7�۰sz�:oQ��w���5����M�5=Z@j����h�4ع7A[�A�Ӻ�����Q�Yq����\l{�s!~-}ƙ��w2I�P�>=�-�0bO�;]�43������,� 3�K�K�غ�rn �X�*��t�� � N��Q�
�%V<��t>�{�e����h�h|�
�:ؓi_7s~<��-�ZuX��p5�n��w�q�TG$�'��)�yq~�k6R�����[V�����a�#Z�s��m��ɜQMk������ŧՙ��-�'%1Mp
f�=���hA}vR�g��޼�G�Hm��2b�8jg�A��UU87E�F���z����FaUI]�F�sW�H����?W����8G�l2��+��|�g�zǙ���b��o�{8o"�������Xaj���-�1��	�|�	0N«��Ui���U��s++߂~FQ�����niR��ղ�#,+zm��O�����##��m8#��o����uD3�t'h�������1#��]���[J�L�� Tv Du.\��^�w��77?�b�LL 7@ٗ����Ik�f)��JM͂)�9E�j|�"��Ld�8T4?RSS�|}�u���TFFf9�5I�Bzd �m.{^ڣ�0	+�3��V�뫟����!�D�bO7ޕb��H[��,s;|a��LSf@�]�X�����'fbE��u_�f���/k�kX�y�[�.�sA�`k�w��X��kN�3/�2c�
�[N��!/�WHw��-z��J7c�[�k�AI��;���]�z���m�lHb�O����3Մ�����)߾��������.쑇���:22�VWW�A��8@��l>��;+FF-K�ڌn�E��ZLT��b��y�~smځ�U���u�����6>j��wP�0 @/�Lo�ײ���$�P�o�c��g�.�]�0���]�Q�\<$�<�B���Y=�[`�^������.�Y�vn�i]	���g>L�=�uQ-�J����!����?fz�ə}�����{7��:��O���sw0��\�ڊ��o�Լ{�յ<y<�e����wp�gZ4�V��\W��#Lm���Q�MU��e�z�8�qK�2�,��!y�#�E�Y��5��U�;���>K���n����m���d�n׺����:�꺛���7�ʦUL�qN������P��`m���~�PSE%���?����ElXx+�n�P�J+��O8��O#_�h��n"��1�~kk9��n`�C�	���74�k�ZUi\���3�K?+������!�`���x�	37QAP��+B�b��~x\��yжͭk}��Cȋ�3��	��A��O=�*��{T_����]j..���X��0�י0Y��0Z�����ᆴ8/�:�ؽ�%����R"&؆Z_՝�OY�v���������� ��*|����f���D��@j7�T�*U4C���#�Ō�׋���둂�x�L�\���ZI�p-���N�Wִ"̞�wrr휰���Qb�6"�L���G���X�W�L,�����Ӧ�F���D���5m*��J'�7�;n�gD�b6������p� ��d����2Q�`q�Q��(�6�f�ʇXI�MXK�$�w>�+���)A���Y�6�}�\�������M�N��c��	�_�jYQ�)m���u��\���w|���l���=;4�-�,���Ka	�N�W�,7���N!��]M�G������jȥ�|���-i,/wQޔ�'�ی�R����~�k�;G��<�r���m�L����u��/��8.YNpn��d��l�9x����+�4��X�G;f;$�@�M4�Z�gY�J��+wܣ�2����Q�u�N��7W.Eǂ����Y��������D�����Z{��K�vw�~i
������f}��ܱkG>EP��w8���C=��D������� g1���z������޽drۇ#��ш������/�:Z��<p`�ҋE���aD 6\����*�������<녽�� ���mF?7/Z�JcRR��u�����n�o<(I���+�񽲄�A�悾�9�[�q�oxؽm���m��gD�F5�'�L�h넙Y
D�4&O�؋���TVs,�q���.���L��?9@�e����9���M��/EJ%g��k<��;���D)�'��U���G���%Uj鹲�q�%����$A���a៑;"���~�]n�RT����ݽ;�p5M��.v��^� JUZV.�C�M��K�<z~E{�r^�THfc�y�񄟃(��!D�[Ib���L���,9i�S��V�n4=I;y���w;�$���{p�s����mpr����}��4�zf��~�a���w��o }��
C��IKy&���S���rE$�G�:�tU����m?��t���O~�F��|:��9���Q%�Hзu=k�G�~Rm�+J���'�h�/Q]MY���H��eG~&��`��"3��f+��|�����8P2���V�Jc�7&�SF�ґt ���_{�8�OM��X�ޤn�|ā<7�P5qӇ�]�]�J�޽^��<I4�6��q�1h��(����*B���D�l��|cOSQ�(��t#0�U��%��>,����Ae#6�@�@^���[(ߝ/�s;��M�����X�a�?�[-6�q
���2�6-��`Ο��k�K�T�h�{e��~���W5$�#��Q�'�[L��<�[�?n8��yUH�lz��e�׼��j�������f�V����,�W��s��v��3��BǣD:��J�����~ml� �������Ϩ�#��3d|	�$I׬2�v�f�P��v��R��T�l(4";;�bW�3�E�/��΅�Q�g��P�;;�x�$.�H�Ծ�B���6@Mb��̨��H���r=:�j���9-5u����;�]�����!P�1];��/�����-+��^G@Eis9�p����>Z(�I���u�*]�+��1��"�B�lw���V�u�̞�w��?t ~��)�)����r�y�:br���|���=P`1�~D�������ߐ`�j+��@���a(�������iP~�bΠ��B��{w�ϓ��� &jjj�X/��X�4S���m<������74�a��,�=�D��0s���ͭ����(�XSG��"��kD1�U+�����,Vz���Wh
O��R�Ú7i�-���K���UcQF���¦�g�ˑ@���MǾ,4��_���;�jΔ�Q��6y��tȥcgB���髪�~���L/��������w��AX����Y�ղ���	~��w����wn���������N�`6[]���Ș��o��Ä�Iד؁)�+���Q("Ӥ��^��v_�geI9�Q�g�a�ٍ�F|�y�u0)τ����v{���	4EJD�P� 	4�N������vC�8\]��N���1��'|SA�n�Ƴ_�/m@�q,܂�\pĴ��-8S�ߞs���M�x&)I(?�\��v�9��_���T�U_NB��9��ɹ��r��1B����ϯ�h!_J PW{p����G(V�3
Ŏl���}EEEq'u�A��f�s P[���k�{�G�<δ+�u6�v�Ⓩ�c�|�ok�����Mh�����T�A�|�7�FuM@H�~�~I��Fk��1�P(11�O��{�t1)i?D����t8���M�ٶ��A�,TW�h�u�w�xI3����W;�H�F��
'��ID��
o�k��@�U�U;Y�@NQ[��<��Dx�|��I�����^㇄s�bϤ�
Wg�~�Ӏ�̫��w�X��y���a!����>�켚ȗ��r��E���[������
�@��C�f���v��TgS�pg�0�r����M�R�������nf�����]��'Ҍ%3Z�t�v`�N^1I�Ήr�a�~b��i����3����r.,�b�ʹB?Hn��p�Q�&}����@ ^�3�71�3�Nd�)�&'��~� ^���w(�<=���$^�A����#�� �")�C�RO���!�х�Y�[F[>�I�mmm>jv@ք7�B=HFs�E}pa@�Q��N�桼��Z����������9�c���ʅ�W�dt'y&�.fO.��+��e��l/<i7YG6u .���m�!��o`]dM�ۨ�譊|�_�����oȸ�666��5٤5�Psj�"[H��ƃ�~o��1�l��-ދx�2�$���{�I�H�y��?��8�&\�!�q�U�f:�Qp}�_6e���t��N�?�]מ@�U��w���¿��8.�\#��:����%�\[���<;�U����k�(��{½�?�6G�{ߧ�ʝ����*]���k��a·��{T�>��f3,�(�5b�^=�R�1:� ��]�!��a��X5�L��Ƕ��g@�Q�քJ���k�I�_��=X���`��Y��L�u��L�[�4���^��BM&��)�����Lq��ھ��H,�+9w�LD˧R��)�S2��yA- 5�i�XBd:L����甎�̨�&T�MkS�zE�j/�jN�閙z���w�JhS�,���y�mm�;���.��W�/�ە����[�qP�W�T������f��`�+�Hw���b��x:�$v��@Md53s-3Qa�|]@���zN)�l�m��Sքnr�;V�H�����گ��s�c��[�V����E�&�"��왤�����~�wAuu�D���3��xD�@�{��;zs9��Ǟ�mئ��\0�=���'��d�w񍏯of�ô9^z����@w�iaouu�3�m9=Xy�ȸ���G�+/�v���3�qU	�a�xz_ �o��B�?�ƭSэ��q�wc�:���x&''��2W\jE��~\c%m���}�i|ڃ����XX�h`�&��C{?�� ��;N���Ng�\SD=�r'!�K�B�FK��{}`���޽�x�q!eW)�2{q�r��)7�!��_�eN`t��9����|F8����C1���G>/�'שXn�Т�����Շ'&���qKyn/)��N�b�����|�͉
�Z��NI�"���ҟ���c}�gb�3��!l#^� 	������=�Ο��~dP��\��JW
+PX����U�~`TX����[_W� 1׋�t
�b' i�ݮ����N��qf�P冀?nV3�#��Ǳ����㻃�*�Xk�>s��~���Y#vʮL8Pa���T>�3��y�3�#�Bѐ�GM�ʖ�񉐮�B6��W+��~7�.�kǀ����9�g�� ����o�h�ŌV����	�Ur;�	},��P�h�3vε'�uԟ��i��f6����*Ë��7�_�~srs��H���?`a1q��D[
�Mm��5)�ޡ��e�lX���j�[��(X�Q�c��(�fhx��
y��l6��w��	�ZW���$jG�W>��j�mUl��rP'��V���Z=?���ib�rv�9����L�����î�p�X�[�[>-�MuX(�x�vZ�H�]견������I����]��X����j���G֯�nI�>��꬗�q� Ɠ��|��g��2d��S�;��6~�ik�ؒ���W�oN��O���
O��pV2�=�Զ)����I^���3�j��d���⻐ٸ��n>X�E���`������{�]W���N!UV�y�Ӆa{�C�:�f#�w��uoee�z"7�^*��J�UƧ�Y)����޲�a̸��BN��P�W[�Z{q��^���$b�6�S^S5�1�x���;�k����������lN�T������]�@�-S�/�5Og&����'Od��m�Ѡ�Zc�@{�ȍ����7_�z��;�E�d���q~�޾R�����3��ȜR����l,q�Y[]��틆4ҚL�rUS;�$���U�������E�P�ʻ,�;v��;{��*N�����>�~�s��|5g|,f8Dx�8W�W�� �7,L�"��[�=�����ޞg�>"����!/����V���m�N(�A��_�������1�JɷWI��0v�\㽊U�^w]&���ݜ��vd���}ON��K���٨s�����^��;�5	��Ѝn�#4�B�z��[�.��zsV�f�˕��ž��6�ψ����D��4mo;HJ��W����2D����5w�P�oJrG]{�?)r,����E"R�wZ�I��1�a%��G�qS^�g��8��E�'F����l�/���$�ú�x�_����yp~�(��I!�4�ۜ��妁J�ni����&L���q�P��ee��=��B�&S�k�sJc֓|��m�2��}�0�nb²���ZL��{[�u���/I�B,pu�VL4,,�wAdm�N[���X�mH��͓8y�
���%C��}��C�;�G>�^>�n��>��֖]���:�sp�%ӗ�*V&���s�Bh�)�6I��3Ǻ�iL�� 58�>m�kFn^dq�b��Vs�
�$������c���:S�|�,	"���囍;y%��%טHY���b�#[��Cn,��ͺ\2�vpzS�2?뙪�1�C�[�V;��/S��x���R�ZЉ��mnג�a��<(�"��?ŝFrD>���T-C�k&�NNN"O�^�ި;�������E�x'�
��z:s����9α�(?w���<|e��Y�R:�]��.b�_,��c�Z��"d��� ��m.(}=��C�P��%�D�í�z��.��w� dկNve�G�������B�� ���C�N�9᝕*�8����h��ְd�����!<6�2�bs6��	�F��>`^æ3����|cc|'l�m�iN��ŨJ��:j�� q0SI1	���po���x�;��Q1�ު�+)���v�;o<_��i~H�Yg��l:��_TT����}�GGG����(����ã#�h�����ݱ�Q[ܝ�+���mrܓ
\��I+<fh�ˇ]N�B�:�7��.��B�&BCC��/�Ϗ����Ȥ!Vr}��z7c4�"�Mo���E3���*@]�`(x�8�b�jX�2'Rٓ�=��#
���$�P�!�C��(�u-��%��pz5+))eWV����,�G��50����mͨ��Ϩ^tsк��)�{�K�2�	V#^�R��<�#���:<̡6�f�*"╚����wF�l�O�`fv�h�Ä�U`�	��wh`�;��=�xSDv��L4��q?Mt����̗b~Ԏ7AY6�Z�*�l�q��43���YTt4��{c1J��	( Pk�® �� ���@�9�L9��d�3i���#NE�99y���fy����mB�~FJ0r������a������;f���r�����*+� c@�{��R�d,8�����"��لV����?S8yB��Hˮy�J ���.�&U[����A��nD��Q��qUe���XUV��M�Yߤ���i��}���i��g�e��敱���\�)	i��ي���F��~8=�٫ܯ22��{��G����k�����Z����RF�Q&��՗�j�	�,wyďp��&S�o���|����
;Zd]}��7���ER��P���[��{d�'�
j8~0��q�5���C���*��G�_�E�}��0 %-ҩ�t�� %�C7��%  --�5� ݍ�� C7ݝ���?�����u�#fΙ��Z׺���^k���H­�T����<0~�{x���]�@��ŀ:I>o����)���ا7PR5�\��
7U��I��@���,��ǜa��C�h�[2wr���D��p��K��R���v�N��T�0/,,������Hq�ii�@�Q(�����to����
9%%6h�e�%	ː�����B�)Jr�^JC�`�1�g���~�W��Yɺ&&y<8$���'����f���X����
MxXeC`��k���Y�0tW�%�1���+l�.U䥦X�J6jW�FyHO�wQ��E����w�N l'$'���V/�y(�Y�,JX�t��g
�$�!���B�Q%`F��/��V�%��_%*�s.��T~��		��Xgk��+~�����C��P9���~P
ʱ�M����I@�a{��+��]!�7?�i�>0/��%�qS�O��ˉ�ց#����45	��MHNV���0� �1O}*�}vy�2J�����`���9�eIB2V��(~y���?b��w��";Q~m�e�CF�y�����D�|���T�c�oS�t��O�L=���/b���S�_�V��� ���{����)9s�P�l�)i�g]��$�?1�in�r��z�;�O�M���/hȎe�NA �*CVe� &T��t,�Ѱ577݈��F4VS奲�Z����ĸ�zR�t/��sF�i������?��/�`�jV~#����(.�a �\��G�|UK)��"U����������f��&��^�%�S����M�V8����d#��O໔���^p���ΕI�dW���[�\Op��%]�R�LR�m���&t����Ñ6�PWb"�Փ�A�z2��]�!���)W��w�f*�\��K�1Sp�׭�&г�@D�[hN^l{������t��U����x]H�t���c��X�~_���:�s�z�������O���([jL0/�����A6�eK�T�¶�e��>)�t��j]���W��S���2EЇ�!G#!�gV��K��	S��5~�3Ss^ַ!�r�5NgX���/-��ﻤV.��U�;A�Y��1q��Z�%��,(�ع0V?̵?��W�	�b��5< �bE��c�U���1j����Gm��y]C}#*[�
������Cʎ�3���d�G��@uܼ�j�
��"�c[��5�hq����͠ә���M�:T�~\��w�W1,�=k=�+�_�v��}UL�D�������d垿;A;��;����`4]�k�����X Rz�~�덈 �[kz��g����޻�d���@�B�굺��j5"�=N7i���4��B��(7[�mS���?�l�����l`�Q�ط#�p�d)�ȏ-������+>�TevQooҜ�u��|�L���ݛH�sy����Hl����M�ꍀ�b�_�<��� �0��wr��T��!խ�*��@8�tw��Ǆc5q�#�`5�� ��� 7�5�m[���4���f��g(��L*-���1{)\�JY��j���W�m�ȕܧ���TJ� N���E�p��(�9�E�]�1�m�t�t]@p����]3�фC���P.�L��x|�6��{�1Ez��%��4�}������1/��u��]>�&YQfI��X2������c}�8�АQQ��DL������6L��)�M[lM+��̽/+�^���^�%���Q#�6�N�f�&�I����"���@K��\O2'?���񡧧ǩ�ގ��Ĵ�r;����KE�������#��;�U7��s�Y�ߏq�f=p?M���Ec퍍{xX�N�X�s�0fwۥnv�"�Km_]�sa�@���?@�1��>&���p'3[4�3���y��R�����aP!�dG8��wyO��ѵ,G$\�{R��b�le���݁��A�����uק~�ֵۤ��X&��'��M}���|3�G�ڔz����wz�x�H�8��g�ٹ�d�����]�D�K�ޞ\(7�����"=/�8�R�t��p�r��e/stX�W����5���/���e��,�����BO��|߆h���/�1��K���Z�^�I$U�z��hɗ�3�d ���i�������D���j���ӛsIC��z��w���EJ��xYا�<}�g�}�.�:��{��^.)]�Vv��2
eNPD^�ߝʑk�!&�=�v�.�`$j
,d���	��Y��	��c���
\���M�߸�ۃ��+�����J[�U��!L���	X��-[�p�sz�%}L0kB���v���&┿�Q�~�����X��L�O�نI�Rz6l�>��U�뇌C��a�$�	��3��3ƊO��`��V�d����5������@��\e�:L$��ޤ1Otݸ%��0�.-"v��^F�l��~u����?��`��rS+O��T��2���
_K@_���c|ȍ[`E8�}�{����ke���˖��˱�_� �D'1�L��
�V�0~y|񳡂���ߒ�+<v������)��\Qf0��ǡ���N?l��6*�yM�wY7�X�?��h��*�:F/���s�����&l�>/ �C������h�ז�!��9˫���Y������>��U#X�P�C'U��q�G��|�V�����U߉w��#�iW�M���p�+Jq �����������C���{���K���ez�-�xq��Q1��#=m0���2NID��vIi���Qb%�]��E=�����F|��[��D��)���i�ɅZ�|��P���te*����F]�]���ϲ=c{@x��Nh�]Hh�lEG���F���]�#��98�L�_}wu#��/�)?/�c�_������ʗ���pq"W���K�����V���嶋k����3;|���W�`}�)�ň���`�gL��UF�� !G09rg~1=��G������ï�>2�R.ے6 o@���_F������%xb��Z��^r!�S��l�`o�.|z����؟�t��l>+Iѯ��R=��d(��s<�Ye>ā�,k$t���\=��E4�b�d(r��w��C^^�h�"px�5Á_���7L!�T���aK��=ж����,�ES��:�$�]�ꪂ��,&t�O�Fk�þ�>�汋�ٞ�;I>��y�'��Jy����j��B�R	X�7M��5��X��OmW���s&�߄��H 9�j���T��W`'��A]��u�OVg�d��"�����Q�*-��"�/Q2�z�1-�H�|t{���y0K�+c�S���qm�N�҅��|c<_�qԼc?y�NW��i��]�ժ��
�k����+�������;���g��^�@&p��c�����s�{t2�$<��V,�����D��lJ6����}������H�1�݋����#�A�p1����L+SS�i��kri���M�����gzZ(����h8�s�����x>����'6_pJ��ZUN������<���#r�Ь2��

�>����0�-F����Pt&���%m�Pvz;u�����4=t/g��݆<� �5fcת��Qh,�3���;nL��D"�O�5mQ=C�G��@����N�7�o�M+�W�|Ky��m+ecso��@}:�H�<H $����21%<��{u�!Q�p18��o�t	'�A����0��p4�ݙM�"��_�*��&��$��Xc}RE���ΧmDʖF��T]ʙ���^���o��)%b,�Z�,�Zk���l ��R)�V��?���.z�������f���閖��[�S*�#b�w�L�������i�rɠ)��c�BI�Cy�S3�2����Ù�q����EϡMe�B���ᒳ���l�6+d�3w∛�:�V��.!�̜)ρ�;fD7��C����^MXI��u
6��k������W��Z�W�,z�d��n���2?��=mC#Q��.���,Ӭ�5���8	'�ɾf�$�l낂=2R�=��<.Z�&j�o��M�ոA���|?,�ߒ�����Er?$�*;Z�m]�l8��nN����nD "7�g�&�L��=5��I�b� x�(�:��� ���Z��J��jDDt��K��L}r�QP~f-^�m/��^?R�뵯���{_v�RA��d�޿��#�����~�P��h��_OGl��ؤ��F���Y�2^	��ń��M�H���\T/�lq��&�V����}xce��&}$d�|�l���g�E4��\�S�oLcXn�$�o|/����L���Q��7f\�;%a4n�+�q���K�(�e�M�䫞��j���,��I�#pZ
�E9����X+z�߰�It�sd�#/����h?ȝ�H�y���M�xA��zU�Y"�jC����>�&'%�ȫ5���൚�*�1�TX���B	�sq�g�
v�(���(4���]m�%s`�M����==�����R��q^ᡭ\�&��B]�w)���-%uc�b�?�2|�GZ&�zIi��у2�N��X���y��Z�U� �Y�ar.�GN퐼V=�����W$cL:�f�Ѱ�o�X�σU48ȥ��l2Ѓ�N$���}u<���!&@y���񚂁�UYW�k�jx�ښ��*��A����K?�Ǖn��F�5�;*�+ĩ�+S�� ���	i�1�ќ�ߚV��3I$ o�n��l�e`��=����p�n5���^�a�l�l�O�eiͬc�E�mW��W��,,5{��Utd
T��Yg���b9�g6����Y��"T[Q���z�q�� ��"�u 36���߿���UUȠ��ݵ
zsT/I���F]ؚ,�#�މ�Z3�W�n���ԣ��c���h����H��R�_���.��b�]da�S�엫���
��k�(�Wcf�vg������ x��ݒ��#�[����� ��|�m��M�vx���hV��N�n�Y۝0»���r�V[ȈvR0�B�w�m�|�����l9S0�]R���+�4��kV�l�6��A!J�_��3w�%a&so�LZ�t����+9U�
u����E�?@�N�����:��DK����:��7ӅQ�*�U2��D���56{*U�lvM�u��V4
�יu?`��͌�)̍�a��<����f7�{�vI@�؜�y�9Re	l�GE<BI2����m�4����C���T��~���V��m4/#� ���m�_��3>����}_G��U�0���ս���u���·0����W)��KKJT��n��Of�k+�f}#�Knl:?r���M_�\�>�˖����%uVW��>���9�R��o|��Q[m�Tu�q�`G>cC0�胩 9��)�v����d����~����05��"�M���ehz�����-����ta���Bۄ�$��������B�:�`�';���Z���X�A�'Ȝy/�h�n�M�R�Y���%N��5�S������,�g���,O�M�w��;��&A�j�S[�:V+xzl1����rXHr=I�/�0��y��az�~��X���q{������ãb`�gj�򉻩���iƤ�R[����&�gπ�f.�AZ��EL��j���<d��	�qK����y.I!~�s���\$ֹ ���.�.���pî5l��R��I�?m�v ��0�x��Kb�.,/�,�*������w��<�ee	�ɂ>A��N�u�i|ԄFTy��1Z�G��*��O��Պ �9��.V��5�j�&m���Cu��n>�DȈ��r�=� �QA�6.�f��+1�������&�橨}~���OԸ��1��������R��5��-��x,?x�tTU��3߼Ѿӯn��z��rr�l=<��F�}/)6��#��H: '�d�~�v�z��$HT6���8Kٮ�M� j����q�$.��dk�^-)��ߨz�ǃ������Q�^��U{:����= ��n73F�(9����\���鲼��"�X�A-6���<B�L+��&?\񽅟s�0�w�~�Y�B�j���jf`P�V
���ܩU���eUK�`�~m?_�QxquV���|�a(�W�)؏7���CE��ې�@?��P�������|9p�
�V ������-OS=�< �Z��ض����X��6|t�(I\G'$���J�շ�:}�$_��!NO+�����;ߤi�� w�;?��U����hE=w�oh4�� �|�Y������/?�,Y�U	�-�z�}�ﷴ�/���ي
�-�Ļ�ECD���e<�~0��a�n�\������ǌx��#A�i4��_�OW�&�md�`ŷ,���3\�I%��??�e9�:8ѝ�9l� ?����^�28�P(ޝ�(�l� �����M���!O6y�E��t�����{���He��Y�{+U���ʥR^^�<�&CØ�5�O���x
M� �A���Ԕ:>��'ild����/n�&@�sw�M�������Б�B�:��J���j�qvDȂs����&K�Ӆ�ʣ0�55�����oomu�%�su!k�m��i?p�^��	�1�$o�N�:F<�\JO��@�ȯ��$6�ڦ�1���dL4��� b���@Y�+��Q/y|wvVG�9���~V��u1��`DKMQܗ�=%����/��a�0N�n{w[{B@s����&�M��'�K"O��||���� x���f�-�+>���oADj�߸.E�pi@�v%	'�0�h|�3�w� �Ns��1ۂ���3�#�3Y9[%k��m0}N�$��zWx<h���]k񍾊W"�P�`�%�R�_8v�%��ѻy@��os�t�M�H�0�j��hm������ m�<�_<GAA=��o�R���ii3m�����.nnOE�����T+��&��Q��;����4|(W�V��P�.cV�&1�9�I���;w0�@�4�:VѪ��QQ�'�O��!m�ˣ��g -wA����7�1L�!�+1�ŀ���/etl��kDH\ �`��p��HP33�bpH.��#��ff�!��P@! �ҁ��4M�놭��1kxpp�q-ZPC���5�8l������~q�_�yϾu=�r�G�ng���e�ۚ��W����q��3��d@��ʺ�w�mie̴f��^�a�q��;w#*�m��YU#~u˵��憐�]&��t�gX8��PՎ�L���b�.=d�#���[����<+km]���tCq9=�h �[Z�L0���ǧ�!}4.r����@�0ԇ���&	A�)���\{hE���%6�6o¾SL{��]��ӷ/��.=�~ZB���g�Q�[�/Y������79'q�홡=a/Ӆ<�d�
4���� W��d���/�9��$��xG�#�	��uܼp�jj�m���00�{ě�
��Q�(kh���*;���x��x��M6'l��������>«��C�t��&���W��t{�
9*eʟ��T��(�[����@��[h��`1�-Ú-=?���P.���9 �{��((���>����|��ܸ���~�jhʼ���5"��/I���1R��(�3(����A�D=\�5t�����io�C������Q�����a�L��P>������Hf�u;_M��L�����F�I�eIQ�"��!f��P��8�Z
�Ae���Q]�����>�7:��A��Y[[wW3{yyWTP	�K<ZF6�{��j�ذFC��Gd����}}p�Z=��υOP���O��mvAT<�f���/��YEzǼĠ�x�9��s�#��i\
}Ryb��Q7��Xv����4������*�ڟu�^�V������Թ5���Mw`�)��ڻ�������B���� �U&np�_��PX�wtw(�O��̖K#+Z_��:�޺2���-�[+VO� ;��NB}(�⽀��Yu��9�2�M���Y���?�u�jG��]:�Ь��"�e�C����ر�J�����-kj%BR���i�4 �p}�_0$WI88m��g�L����'}/��{�f���`ͦ}�Ƚ��_�EA���nc�n��z��W8�%jZI�����Ǖ9��������S~������nc���e1ZR�����
�"��-2=C������+Y�Q(0��v�7��a�ݚ1/ɘ�m���b�{�t���T���Ȼ��*>��
��ك��.��v608ג�L+^v����}y��s$n���ϑ�����O����H�Ѧ���G^ݒ��T�����B<h����$;�!��db�m=��闺����Y�I�b�Va�-0d|��oW�Z^�cV�Zpe�3��5|O�˰7W3;;;���8�S��bY#p�[ҋ�M�#���h�k����X:���'�D�e5��}����ы l�c.����\ ,�ՠzfχKL��僾پ�'�	�����B{?ۭMe&���.��αb;ww*2?a�⁪FUsK�&e����A-ϫ��@���ps} x2#|_(����A�D�����6V�N���y��V�e�񠗋��H[��&u���	��ݔ3�:���D�}���	Ew��Zkh�pQBr�O �+f$4>�򞧙��Ƞ��=�mگ��
�x^��}�Li��5Ϟ������ۭ{���6
�]������2Q7�T����}dRҀ�Gt��@8n�d��z-�jÕ��3l����p�<�M*g�j�<�6�h��>�h;Wg[*��[
X@�rr^zqc)F8T�մ�W�l��Bt�Z���`���l?T�������a�������1b�\k�9���:U�.���v��ݔ�/�k�U�G�5�,��
ӏ�+�_~�g2��0��Z:0//褚9dK�r�Г�P��m��*��S���ۥ�wOe�R/��^��������y:cp�g`M�s�G� J�+��[{{�W�ke�Gp����d�s|h��]�E��(#Q��uuu�?-�����������0�+�dM�/�Ua���~?[��3���=J>��4V���Â2�W���.�qJ �mW-�����k���Ʈ����H�w#	����\O�բ���aX�)�9>s�Wb����-$�g7ڒ�2�������yb�=�a��O4�ZC��6���ióz,�X>�V�*�)�v�7x��2���6��q�}c�5��1���.�s�8���?�s�.�A5�^�[�z�CtZX�/�X&MoR8ZZZu�MB]�J� ���ڳ�˟�����#bp��
�;�GG2��J<�V*��=^أ[)�m:�����.^�2��kn{��i'YЪ�ϐ���5m�� �2���HK]�2�$�p����Ns����g��kb�I��\����6���v諱:�w�x}_��{z�z���a"rs��q��z��~���*�^�so�l��?��r�?��s��?J��΂��P�3>�	p4��7p�,�?V�f~2�ݟKC�"��TV�2�}yu���7RX�&�]�?8+�}��F'D���[����o���P�Y=TL���I�3
׫���[�ĵC�5�-��@�к_�Y99����ZVMwU^��^�ék��O���0�K�|���pՏ�ɼl��:���i/���]=�'�_}~#r�.�g������+�EoW+�v?YY��Wz iV��
�ޔ!_{���������cQ��^��������Sn~�e	����9�O�w�p�)}�����޺l�����(���!c"�jN���hi{����b��M!+^�;)ӽ%��>3�Ĕ2o]���"�����^�,Ȳ��s��갵~�'A;���K�v���%�V�>�+���v���m�q+\��H>^��\g���a����i�7��������$�0�� {C)��{p�;k�(t�g]l�Ũ��sK����s%%%+�b�}��t�OtB]]]Y�㖽,�d�0L�1�=KI%0�$�~0y�3�mI#��T��&���V�����ɰ�ӽI�u�۞x�u7�����^�o�Zb������
R�FQ�s^:�y��0����<&�M1�"��+܆Ys� ̫ ������k�:r��������ܠ��2σ��S��r �����/�q�A�����@�����6�X�����D�b���y��- 'h�痗l�^��9��h[�w.���tF�����"c���1?�B�}}%BC���;G ��Y��-�zN~7,��'�u��:�ҡ�6q��0����5����(�,���9�L�}�{�������#5MEN�D�s�T�������0mz:<Fh��63m�@;P�E�Λ�QhT�.��# �P߭���!!!�1��0�ӥ%X����(��g��q�h������2c"�l�U"IȯtɃ�ɬ%�n}��j}[�(ւkĄZ"�����%
J������$'&rp�K�vL�I�Ku��"��� ؘQQ�R����U�6J��v�'���Li6%��>Y'��&���q#|�M��W���{�����3�ǥ�/�����}��%vh7�j����� �20P�&1�KBf�l�c��b$v>-l���)//���/�'��>K��ٻ�*�?u�OS�90�Im�&3�BM{jH�z������FM]�9f�0W�߬�IцY�|>���g,#������cT;r�]T�9U���?XЭ������GF���6@�� P	LE������?lW�����閪��]h��(�a�3g�t�����<(�������b{f{?L�r(�6���%eN��V�W8��#)h��98;e�Ѷ=�k�熱?��S��Q�'��� ��x���<��[b�����'��M������og�M#��%�/�V�파^V�d�����G!d�@,�$j��)]��Vn"�C��dhE�Ϧ�F>��{�S�x�Ռ@\�'����N��M��D�-�l��34�d�$`��7b�o�l��Ox�e�)�۝�����a�����/¬5qR0 ���=EL(�QzPZ/�iC�Li����1<]B��?gm�C?DLwx��hn+g�C>��߼��<?]��������ic	�������\�&e�s��i�����罹��S�p�gA�8�<V
F}8Sb����p�Vȫ����ج&����-�&%�ɅΛ[�f@�P[�`b��
�>^�g�����xB�l��Z�k�#S:t6+�4!Qi:�:��֜G����E���`{P��I�nv~�uT�"����=���N-�`;���Y>�B���&I��!֤��������
��llsG%�V��MV�0֨@R:��-w�>:ĸ�VL%���]fA0��Oj���Ms@�U!e]�k� ����������X�V���V7��O؅�?�@M�x�%5�[j`�ԋ��[U��'9���)=y3�>J�B-���-`�N��)j�Y��NI�p'	�)mr0��YU��o⅍�~w񊬮� \��Zg�ʟ�,�o��5��zg�����w���[)ڦ��}�@E��}�m���ӿ�E.0�~�-��>����@��m@+/����#�������FvjL��k����ܶg#���6Ƌ�/ʸv�� ܲ�5��edЂ����������u|�ii��L�>��M��L�^ե���A�*������j��u���G��^�뇥]���*��-��O��<�/����sQ�MML(��v]]��"3��N�@ ����6���5x����2�̥0����I$�h����ب��Pǚ��""DFE)X|���ƱbTT�Sw];d��7孼~��t�Й�����џ�
�!.A/~=2c,�k���8��!����{����N7%^�7n9���x\��=&x骏/���Hf!�s�Ģ��q�Z]Ѽ����c���-S�z��4 ��S�	���O'�m�����6�|���*[��ʩ�G�����ӧ	�����}���J�YF��S��gT�	����6g��Yi���hۼ�C�cz�@� �,��=-�����0��{l�$��,b}V��p���Q����I�P(d6�ʕ��j�E��������Ԕ�E��&v����P�ve��L`�e�ɡ����Rؒp��A~����W��u�F⥴(�V"##��E�~�A���ݗ�e�����`!��)�y���%���O�VM4鐮��_���OX�ee���7����K:���+°�J͖`Ł��}�����Yr�@��讎�)���[ۏ�#���c��g�3������wY����_��Hf�ݚȰ���K�o��7��1�ǌjJ�[j�s�V��8_�l��s���M�TN�}N6�ᵵe�~�@���?g���uf�ce?9��EKɲcȿUeU�ꠂ������߅���}b�ԢZ���\Zr8���t ��3���Ǘ����u=��.�(�7y����BeotH�)BM��$��O_4�LNL���7�|�;����#�yy��we�c[-��L��ݝM�_����K@=���v'���ht�z���E����� n�A�/��dS��s)X�	d<�ȱd�,��GD5�z��/��4w�j]{q�s0�<D�/פ٤9��#��lT���{�n�����eذ���(�y��-/i�",��g�V5�����@6)�Q�V(k��:���+�/#�� ����*u������I �7���n{��O�,lx��Ř�
>>>iS����nc@)�t�e0��l����c���1�1u�� ����̪����Xue����m���Q��>���⨖5C��ȇ�K,W��V����������d|w�|���1j4�?2�B�\x*i*��1�M������j�FN���%���z �f��qф�_���ڽ�h$	�Ǆ#���b�wy%�n�����^9����fШ��D��6�0Ħ�f9?}�*i�xUk)w%J�WDTxhU��Xiv>~n��ŉ�mR�����r�zV[j�����wo0���HX*#M�׬Ʒ�I)qj7>�+�o��ӎ�F��pk���SB��+G�TdX�����Tݚ�x��X>aN23l������;�����_?�Y����ŀp�-,���$�I��Js�Q{[}�(�Fy�M�0������zt��X��|�0C[I���}w�ز�Q�B�+nv{oi#�y��k��}:����?�I9WR`�����5.�iW�GȔ�I�N����<��~!�a	��Jo�	��/Z�c�m|��p��V��٤; ����Z]'���ׯ�Q#0ݓn�rE%%l�*���i-D��8/]�'R)�>8����ӡ)� c���C8���b�Etm}]Q>f"R���L@i�&�f��M� �@�zf~�؟	���{���_��4�\���_Ĥ���jz����GL�!fk��t~��8��q�^�q����Nɴ/�ə��\\�77�)��5EL����Ϝm��q?eV�j��.��n���Ί�|P��n�	S@>k�w��������fC�wo7\h�PV��/le_e�����Ǔ]��\��N��b��x���+�d��ab��c<d�4G=�FU����ݳ`.�acy������t���V�)�b��+�������de�q�R0ꇹ_�������$�t3m��~�������W~k|˾����
��v^
o�U�F"�V�	"�m��Փz�M�)���i2~]���Q��Z鍭(r�W\��{_0Q�ąZ�(f
=�f7J�NF�]�Ș�@��U�������e�����g�H��ur{ODI��BL��+��+n��<�����S $�F #���q(jΉ�"&���co������d"()S�Uq�c-J�@�6ߓZ�Y4��L�߾i��Ȧ�-��P��a]�=|�����eG��ln��P�Av�c���K���:b)fޟ뮒��I�ZN��@�H-��z�J��W��ʗ�p������4ʎc¶ ]����+�P����p�ߩ�D��'�w5�P���M��_�����ò��W �?�R�CD�$�H&v��[�q�ź�*Zю�`�be���gt�#�X�9X��pw}�bx�K}����/�&ϤR=������|�Xe�ݿ�6��>����̅*���_2�Y䱵~�B��Xݛ)i�M}& ��8F��g����te+�73�mg����x8\B��Ҽg��~8;u��A�d����� �LT�T&�"�FQ��Z�h �k6�����o4�?D�i�:0Q�īA��*��J��ku}�;s�,]�ͨ_Y/�V=6�t�j����0�P��s�fS��Vbw3����h3��	_��5�z}3QrA������0l����jp��@S�>�����k4{����w��6�4 ���n�n)+c���d&�{A��lĵ����1��:,��:*�W)]��'���BA �ҟ����������uL�E�y�
����T������ڌEV���V���upé���1�o�95�tl��_�ϻ�x:u����{õL�1�gX��%���-'���=��:j�p���;"t���B���R1euw�$URI��g�J�E���̭*�ے5c2y0��R�.lBP�ȫUN����ʪ-��N�<C��b��t�����V�C�`�l��B������ �u�4-5ƈ�ꛭ��lM�� �d�����y���ݱ�4N;h�Ů��������c�m�gef�g���%l�FlX�-w'�L��h��w�X76.oﮎ�!s�������8�N�9J���ڊ���NŲ)c�W�.�3��pzʒi"|��'n�Y';F��������v��6A��*��a��s2,���K����Q�yL����	G�M�ػ��e���4�!v�'��P?�����Za���b��
�޶�WTS��7H�=1ٌ��G� Qz�̾�}[�c�D�T��d|�uE�Ձ�/HE�<��U�]0�	9����oC�8������i�J�:V\r+^7k#P��o�g����{���h$�đ؂��W�XX��`�y᧾(E�g��	�)x��|%��Fm�,��s<���R�oqEŰ{���RT���5~��Q���_�;{��3=��˥��Z����X�2𠗙�A����mC%�ʫ�ܡ\,/��\�y;�nE��S�O��x[�����9�Ҽ}�����k��	h���u������������. ����`�G)����@�9S��P�5�PB_�����ͧ�0��/��0��xe4�yirfBk���Ͽ熁�i��Cfkk���*���P��L������&��{���y��{�f���3~�s����`����<mG���[H��xn1:9Z��U��|�ˡ��kV|8vN���#]�
ZI��1��}�KQ᛭ob��/�>:Ff�v���QSĈ�!� K�(Ƥ�KP�F��*�!�^�ww��w�2��(3R��!�$רcDm���a"Y*�(��f~;�4n���Q�+����QS�o��"066��n� �����Wf��O�������g�"�؊9G�y����H^[Z��n�%	�A���E����윜�{A6�RCbc_ �����g�A۠�]����*�v]�Z���t����-HwIs�1z�~��_��Y)�'����*,*��<H��	��I�O:%��q+����h���<C\�F�t��zA��e
ߩ����9����F#�<�fm<����X�� ��y���{Q�� ~_e�0;���c�����>��
Y/��~s�>r'��*z|�e����mz���I�U��'��_�mM2O1������������lSo��~zO�"ŌΤ$�	>�
xIv�.b���\S�㐰x�O���~���6��)��� �W10����V/;5r��DI� .�P���4F2��uҢךvAk��￩>J����w���͖�����@��f����zQ+��P]Z��Q<"]6#SĐ����""lmmI�)��y�ʷ(6����� d�"�B���~���.�������>r\Y��Ô_2�Z��2/����˒z�x3b333&� 3�%�

������dn�׭ �=�>��r��ty�=v��>�Z]���&�=h^i�4��s�<H�^� �~+ɳvٽ��e^oA~�b������Vd�΂�`em���<�0���(�����u愅�yP�U�)����YnY�����Q��_4�"�6L^.���=3���ߤ�����P࢑( G�[M�TBX��Ms��R:��	_]�d4��9_}��	�WCQ1R㧢�U5%BF����v���j���S:-�k�UURgF����ag�ME����N�gͱ帏���H�ښ	O�>����D�Fq���!h�H���:�IF*��	�>�Օ:E>���\W�U8�v�f���`��B��b�c@�b͟����Z$KH�=��2(=o,�H��C�Fժ��c����L�����C��� ��,�B������7��FVV$�������,��,�!q�ʐ���Q�5{��}Z0��;F!;����s1D ʴ��T���������W1h_�m	}����ؽV�_��:����Y�W�ml0\]]��I���V��Td�������M(���^{�{�v�z��w~"�%D�MBB���Y�3S�Zh���=`է��&����h�M�ӷ�#b��"-�t�����XX�D�٭�L�LK3 ���G'��LE��"��v�n���oo�,f��w�H{&�վ�I��I������`�o�]�G�<͇��a��[ |<D:���ۉr�{��~1��8{����mx膡A�P��;����Q���A	i���)A�n�⽠����k}����X�ν眽����}Δ��$"]d{�y������$XyB��H�4�:7%���PtI0 K�&!<$���ȡ����*የY�z��']߷��:���&ێ?� �,������^�t�eĄQa�����:?�$�A(��3}p6���L��$�P˾
���=W��ݟ@��P:PQ�W���*��+�S / |EEE��װ�����D�[�����w��M,O��Wx�����@� d*Z2��ghk)�+����k}��ᐌE _�X���!�� ��#(�3�C
o�h�B��vZ��C� �g�������Р#�0�61��`.����z�ڂ�QUs�UC�T| ���_G�N��q��:�*�P�8SI- K��ѵ�aO�~:7�K��9_�f�+�H�	Eqqqf~T�����X0	�^9�������|֟Qp�f��iM���;�<re�����`����!����4g4���ܞ+S$�pա��4� �
�4�k$�6.�a0�Ia��sZC��_�7����5��F����n��������U����ђDI���*���I5%%��������&�S3�}j��+��(�d�8�;�~�,�<��3���2k�ë�[ퟏn����f�BC��� H��dʤ����H�_�.(,|���+��A�7J�Z���/G�}����CR؍B%I��'����W�v��HGsh�/'JC�������T`=ַ#.�o�v=�L�l���J���KqYY9�a�����oI�4YEE�			@�M>��c� �T���q�gPc?5�� )��N�~�b̭2�}�����X5�@Xm��#VJY��e՞q�d���I5��$:||�B,� �l� ��n��ac�`yw
�����b�������qA���l��	������G�e{D�Jd�a_�*0��P$����4j%�ܩϡ�I�(=N��/����YB��0�@��k�Pc T�^*{k:�u�����#�ƼQo��k�T#���ƚ�ph��81�G>�"���D�aC������+��m�t��f�F�/�d�
+��M�i�5 (Qibc-�pA��@��wN�����Ԛ�ಠKq��(1��������q'�0K�jI�j!4�b����@�}�#,��M5��\�z!��r��ՁF��L��R��j��r���	Z��4V�Y�R�՝8��!�3276������	�D�S^��d�x����nxH5}��hrC_�?�޿�`0����B�-B�xӯ�"��,l\ݜ��n�,���4���nl���ݤ����?%�hd}y�a�
P���'p��`U�9b4W@|lK��}p��X�w5)~�/*�kc5�"h�ރ�%khE��1=����mxh�u���$�]���;���E���~�nK���u��?�L��%鳤6�B(�;���1_��g��y�m��&�:U�*�(�Y�"�Z S��[�3�:�s� ��L��F[˄���Mf���*LXjEV�Q��"~�6�����<��T�ɗJZ9�]�< e�ϕ�)H�d���$��P&��H>�骞��n��~���N ����@���?Yuu]un��a|�XC;�nmz^�m�1�����{���-���� ��L�'���W�ոY�C�~���ϩ�A��x�4`z ��+��@�f+����*��W<�,��3}:Mv7�S5�<��q��'�Շ�S7��g#�jDF����0(����}�j:�l���D��y���>U���a�b@�p6��s�w.����ɕmڡHMeO��3'��%��W|��p�48��6�l@��A���L�B��J~5A
���(�IΟ�QC<_��&�x��b��Zff,��=���X�^.^��W1��n`+M;�����8����) �I���
�L?������3�յ3��""-&�L����pMi�@6S5������¸Q�#�a��R2�����؆mG�ݸ��R�[d�&(���ߥ�Z�q`|������9��˗�~��` �D4ej��L�Kx��A���T���#r�.�'y�aoA�G�v{g��������WNt��_���54��d���O���(�:?*~@~��r~�������$���NT!D�����Cذx��4����p9�	]��(�����'�T��{	�3�{EBN�ݻw�h���Ũ��t�����J&�ݵߒ�.!�j�@�`O!���Tp��=�i�_��i��7޿F��Y�@+���"Ī/w��9�tآ�����NbԶR��مٌQ�����-q��R|�;x�W�J���{���/�_�J��(z��
O\v���N���^JQ�VlՓX	��U���{^�?��Xl�����˜��Ԭ�JE3�ג���8�U�=k����L��V7����k�O46�4�2{��R�)���[�_�8q�`)l#�ga�l�u����Q���@`�s��tᓭ���x��1��Pܭ��C����l��7"�N*v��^K�r"�&-��z�����oOđ@i��۪/��OE%z�1�ʫ�����J�	Ds�]Q'�*TJ>M	��{�g�����4!q���k�q_q<-1]�H��K�.;���������#�$x�)p.�|�yQ����k�@JPvɶ���|�,�}�1R(�a�#U��5���O�`s�ӒXOy��{X~H�6k�_�	tb~)���:g��5���E�H�G��$P�?��ό��&\ɱ��r>1�=�.�=��w���v�OX�7Du����"hXo����UVM�d?4��}W������q��~a7�h2_I\(��ą�E?_ne�$��E����`]�ʛ���ۍTs��4��* T��j�5~ �{��l�/7��-���p&n�����?B�t��ρ8}v��!4،�	��n�����	����wp�fR$!5�=f�`|oo�"��z��V� �9�K�ͼs-���En��w��*|E�'�yaq�&*xO�>�t�x�����6&���O4�cN
Ր���ҿ������������#u�
�:2��	�����|���z�x�gr�lf��Eo�wze���5?���/E/��y}�2�5��__��I(L%�G$a������4��f9�Z֋W��˒Y)m�!6��U�-�E�'�u�	V��!�*��3�s{��.5�����ՙ��o��'�V\���^dӼ���I��F���&�n,�����p�j���I�7L`�*-lcc`�$xs�"�������_�7��^�z�������0<��8#�����!�A����Z���GT{��!5=&�RI�I����ъ}�}?z��,��|>���N�n�bw���DY<��fr&/>��*���1����ƅ��dC��L��0,������(2

%x���T��b!��u͌���
����D�<�EEqZ!A����d[��]��Qn����f:$���AdI��¯��p@��K�<�&
:fGk��VZ�tCr&��Ծ��<}��������/��D�a7E�d��`+++����{�-}X� $��`��qnnn���KKC�,�?fq~��z�M���U�x���/�|�lA���V&�|�4��IH>| ����S�و��s�8��(�b���&''IWS�##�K|V�ʈ�$i�L���P���y���ޅ���C� ��8�݌Ȑ�p{��y����F�7, �����������3/��2���{$��K���f����;<�?n*��p��i����6][��u�͘H5.1𦶿O"����!��}�b�n������P�)��A0���l���V�D�b�����ggS��8Է�B����,)��i��H�]���:�����ΒrҌ���ps⿽(Xqf�cWj\x��σ��*\���Y�FYz�os���1 aa猤���7��,����	x��j��=ܦ��_�'%dӎ�W�Jo��e{�	��r֞l�©b.�{+[JKa����?/����d�!����㻮J��myV ��;�.T��V�owbd��_����؉{_CD3j�\`�����	7��ۧ���+�>>�VV�^�z�ރ+�?<l�SŢs_�z��_DKM�k��O���V��D���&g�b@�N,,|��ΖJ������~�gbn.�^ :/�I8T{+�� 2�����#`Vۿ����Ӄ���������������z��i"^!	��vAs�71�����&��¦Ǐ�u�s��'-d��b�G���n�h������������������j��J�x'������hM@r^D[����F�t0H..���D2�\_z�}þ�/)����s�ks�)�����[�7Z�ё���������6 �.���oM3��&|#�_Y[c������2�03W��ρk�p������76Dly����ŤK����𻻕J��
xg�b�ԁ_*)''�vnWPT���9��z�7g��QzO��S��<57�/9�DE9���e��c���8�5�y��x�*4Ţ����X�5���R�<�9���+&��[�n����G6���8ju$,h��2��f�6J�բ4^��j�2g���f0�Y������~�Ow5�SSSD�2�|� �QML��莃`�(�aT?��߸�͗�BG,�-�CC/��b��]�[[)���~g$��o��}෿���#�]+�j��aؐ�i=�ۙ�	�
\�Ƞ�sd�c��@����3`�K�\(D=��b�B�"�mme��X�gE����V� ���		ik_�Ύ#�s����.��Èm=iS0
ٸ"!���M̡����3�{L�P��w��%qCB|333�F={
�����$�AK�=��u�j�,Tm��A�JL e��sw�<�J/_�zz6�玣��U���Vjg+2Yď�m��ӟ�l���%+��Ҳ999!��ڬ��<X������>�'Ӌ�AC/}�.6���ģ�<u������{2�������{��O�#��|p_��tn���o���8�bI������ǵTY;�1��9���~E*[Q����z�Άř\�V�`���^��:X]��@�*-�}�����)%����d�դ���o�����=녩��#������m�v桲���[!=vXU�*�tj��Ϩͅٽ�k�f�|�'���d�[r����^f�'��ۃ�ϧ]���{�ڣ�?�,��b��3r�ޡ�z�wq�=�����L��� `�ÄiW��[����I�s��lisQW줃F���$���������a���/��-9�R��/����G�fY<z�ڽ��z"�5�g��C
�������Ĝl������Q���x�����/�6�Û���C'#����a1� �R�����5��w���,��?�dpPBBBβG�2� �����	0��6�p,7L**���oؐ|�s$4��z�[��<T��+�]�~=C��Ѵ�� <�ө��ℌ��1��m-D�r\b���0"���V^����
���!��� �����?H2j�LL��J$ڀ#w�h�A�zt������rtll7'6Itu��Ve_�Z��?e�e�bh�,5�$ꎟr�!��t��\?�$�ﻻ[�������ĥ����C?��u@���q�*E8��X��P��k��sM��H$j0U!En�ͩ�P3��VYI�~{zʳ��M������o�l�c)v�m�8�۞�27�˛��bw�x�"|W]X[�;�5��g�3X��8m����;�9�Lx+��e�F�b�;�ukp�����P.�.y�4�XsR�j�k2�(�	�+�LL�s�Q�����Xy�͠`����D�@�j8PaV�f�o���_���y�zLa!�� ��ag�{�il�n(����G�{6
��؝_U���7���7�M����MC�5���E(ΦD�i�돍5]Z�������	��v���=X��ja̝e��wQ���=&�=����U�F��2D�~��;��B��螫�iZA�.U_�iˊ}6�@��Y���l ~r�wV2��JJ�y_4˟��m;{������W�m�Z�����^����?��%��e_au繯8j��� 6��F
����h�Yh"흡tD��s��pgt+m=W˗Z�Xn����̥V��\4��'Y����֮2���Ƶ�38l��/��x�*A4/������xI�Z����=� Bڼ�g�.-��VE�1%ORCC ]Ž�
�sx�"Câ��u�y�)�l��c2mX�c �( �"����ޥ�� �4.k�_�T��%�'m{�L�ў�tNn���D�` �a � S]� �q��~�9�H��6_ϊ��?�>��&�B�)gt�c�����
#��R�$t�Y")q�2�8}P&Uu�*Vi"�����=���U�	m�����B�c(N�2+?�4ΜȠ�*��uF�?{b�
�+��F:_��߷0c��ٟ�?Kk+X9"H�S�����p%��|�#2�h,M6�4�XB]�c��p�b�I"w�G��r�x>�$�0����C�o�U "x���� f�*>�]_'�BC5Nyp�
+�!/�47�e�y'���o�����iƚ���;*��������Xm3�zu�j'�>s6�|�����dE�e5i�]�,Eo/heT�X}%�We�АEз��M��489�|~��<�R^MHӱo߱b�g�7$G����x�7DW�����N����������t%���p,E��Җ���5��ȇ Bq��E�^��n�������߼ $��k� ��`�&1�q*9*9�в@-�d55a����k"ഏ����5��+�Z=+����B�1��k��womm][e�2��6��r�%nV�h�H� �۰���fR�������N����T<�{�"��>�Y��]�*�Z^^�Ũ^����Ҭ$A�����fIxB�j)�ZG���|��Uqz�G��� ����Ǳ˰��R��ٙ*
 V-8�6��44V�<� Y���������� �{�ce��wm}0���ݝ��k���� ί��jN舸�B�ee�z��f#�%�y�w~66l�{sh׫�(�b�v	M47��B���t���r*?����8X�~�~�W�����\��`���B�K?����MѨ��*h���;Qˌ3���ii��ݩ3�eN����t qrz��}��,C���9���L������5:4�M7�� >JY��q4y�$H�[S[�][K�୽=���F�R�~�At�������J����4/*
��Y�[^T�9Wo'ggg����+�f?�˪�į�[�1��\mۤj8h|�s2�{pQ%$v|:)�h������A:�����w��ݍfd�7�h3Z�ouF��� t�d�jDZ"���:9���g�'*q�^�;������U�Y�������)(�L�K�X\��0��OIy���e��L���.�@`ng%c#M���t�;����TW��W�3��Ki`�ց<�2i{�nCCCY;WE)�0�0>��1�g�	���ԵY����9<L٦��~+�C� ��9NZ�;0R�f�>ʹ�h��ݞ�\���ʫͷ}�������i__���C:�� ��'��M]Z�+MJ������J�]��l!.;0[t{�`�sx����u?�{�
�"z]����?P��m⳱y�3�\D��j���6G�+. }˿h/jແ^R�/��NǑm�
�۹i�d��w_�0��}�����LתM���S\��񔲣���9^�M��z�^�c�l�-le�H����/�Нv�r�c�w�n�'r�`;|:��T�n�)�&���v��_O4���D�E���;T@m�e��zҌ����7բ��4^�V�V*|���%Iْ�M�ٯ��(��©����-����*j�ni���7��?�GM- ��]"�l�{��h�ȈU�ƃ�y���a�����|�I�11z̵mw���ƙo��sa���U~��i>�m}/3�z����b�;j����~�����(�����T�1�/�7鐤�<uݝ�{��AU]'X_9}4��~��ָe#T�k ��L��rȻ�����2@����Y;B���`�[�����m�����h��3����γ�r@���s��tF����yX�����봕[]���>�j;�u��̣��涿r�6��}�<YkZI�vwsP��U�s�7�!��[ʀbl"��R��CI�ss� -@��:'�I3T�щ��_H�3���S�Q*�u|şՓg��n�"�_��I�X��Ij�n�#e�����v~����~��¾^&��[}SI@���������ɣ�E�&?��&��^y�
X|��8m��3�,��?�>1����)���⾀r��S�a���펐�ͬ����D�G���:�/�&DG����E?q˻���Q���<������o]��x�XxRG��9.��=Go�����gs���`N�A������1s��kSӣ�����m)�S�����M+����^��8��:����4('bxU�ғD�>�@��Ӑa�4�ӥ|Rk�+.�<�R�v����M�5�tC����7��QI.AiQ��԰�7���g��-�╲���/l@�s��:н���f�rt� ԰`{�1{�f� ��N$��j+�*/�WX����woT�(����	1~ս����,��+=IJ .V��bO�
å�ګ_�aӭ���A\�I��s���(Ҁ��7wR?�̰jp�6����66NV湰�3}9��nWͷѳF���./XZ�	��R�LI>��R�������R��7c�
�m%_78��#I�+�.l�'�9���]���.z������:W

�" �Yl*C0h��=�>*h���v	Kq#9`F�u��ZS341��z�Mtm��(�T�:�3"� �ɹ�������]�N�S	���T��[-�����/ߜ�I35�ȉ-۞W�y��W�*_��41����N~���h��p]�F�}}���wRoXw�ϟ� ��X�&E���G� ֓�ANk�[S�����A�C�e��o��ٹ�H�ă�O2���@dG�6�8��DFtż��5gW�_�m(�^��������P{6����9�i7��v_c?��7PV�N���u��;�yG�z�,>����7'#O�vAb�q��O)]l]���sB*O'��Hx�����|����Nn,�L�A	 ��},*"�doA���i4�����ǅ/���)���ԯ~�䓠����o	��gʜ6n~��=(WhU����	��N��G�Y���q(_�b:��:��b����aaa��KC��
-[��Uh(��?�(#pJ��
s�,2불��V�qVW/iakpN��Hn�'�_�Fm�Ӈ�J��V���s`n��Ҿ��\FThq��M%���UX$i8���JD�V̚�13�sA��R��?rm���M�N0zy~�ޢ���De��vz��/zsϻ-ᘅ�~ݸ�
yxoE��,�HD�L��&D]uK����h�th����G����ţce�VJ J����A�.Ha.�y�%Wb�U�;B�V[�4/,--91 �zǳ^�l?�W���R��`��'�������_�p��B��^�i-��=�~�И/��E+t��1��[����ɥK�ӈ^�/�+ Y99'�%�O��'s��d�ן�"#1�w~�P^���md������<.�o#F�qS�
��M�g�}X�����Fz���m�7��l|��".̦��cΦ���n�h_��j����}�,���ѡd�,�]%U����^I5,+�;#m?���������3�f[O��=��ӧN�cR�2_���p�����UU\���:_ �#�@.**zN�n@0��Z(�8�������@������7��	m����ر�O�&bb,$�qf��[7�k<ql��Ǐ���6Vι�{�t���ﴝ����!�8M��.�I_�f"G�P%�'&�8X���t���he9~D�|�5�����Db�{�����T7`�B6�4�A�3rm��|����Q�Au�ĄN�%B�<��,�D�j���N�I64>���r]�V�F����i����)r�O�Ǽ���G�ůiC�b��pQz�*݌�al~����e�����X��v��޵�O�>��f�^��IO�E���\��{� �����@X7�s�1��]��z"dg,bty�y�\If��K8nu���6�M}]�� �]��ȑ}Qj'���!ic#3,'����e��ER.ӿ&���9�ǫ���Տ��~5Q�,2Zb�:�Ҋ�f�mTWe�]x)�<�����a�n]�~w�M+t�j�{�(s�����~�k�!',��?H��cC}������(J�'�߶$�ԣP�¾����������j	Ϯ�Lyx[�:���\�$��>5(�U�F ������_�Qo~�7#��Cu��<�.,,�#���5���cq��<C�o��N�@�ME����E�%*<���0	;ڰ����\kZ� �ib��㉼� <�+LM�7�!Gqn�C}lq���t�|��+ڲ���8)��+��:�@��L�
�wz3A<���:1~���]��)��¤u�����wa�S�b��D��l��_SN{��m]��4���AB�Ǉ�	ᅬʂ�������s�\7L����|e��TUK�@��ξ�i����ÎQJ�(��ޏ�ߪ2Nt�o�37
�$ʊ�N~�Vc�_]
��������2e#�/�]ἰ��'�a��R�#_���]��#��ǱqO��G�����J <�F�4v������e�k�.�19�Mơ�証o;�����(��~3��Z젎M�Qu��fv�@;��
|��G葸{���R����LF:�hS{s���H�t����O}����۰�"�'��s~�BXX)�u�S���.��R�;�&t+l��xNp�M���"''�=<Pq�r]��{���ۗx�渺7���(��1��-���;�w�(Ǌan_�����N��P@d�<--3T4gI���Ηj81Ҥ����fؗ�3�|F_o�q!��ߤ�VRV�tL�Q��',��|onnB�i7�}�����7��`�56�C}/�V�����6%H�Y�>�N�>G2�Բ;Gkd7S���^��T��Lwr�pR?����|4i��"�MDmɉ&�.������6��C1�G
p9v٩����32d�NR���%���~���Y5�'7Y���E�L-$He�(�>� �q�����1,��l������L�ɖ�������L}��$�W�UF%�x��`�x������ǽ��GEs�<��Zs��l^8��0Y�����. �b�o�Odթ��.��G�uU�<�w�W��N��rK�|e�&���x&hxt��'�mǘ&h��'��`V�����/b����f�Q��5����K>M�ԛ"*QV��Swe�-~	���g�Ay�3P�3�7�����Tp�\,��(W�c�����n{�J�A�po2*����l�U��Ls��zQ%(�\\���^��ke�~�H5��
����Z+s�e��W,�Ȣ3?P�4~��db�F��A'm@n黼\w�h����c�KP��~S=Q�pώ�W < ��8S?�W27�evka�r~�o�?�x7L��ϸuvv&��l��9(:rde���~)x-Fa���x������?I��7"���U�����x������qg�^�tYi�M��r���A3����N�m��P�OAs�]�nU\gG]��Cf8,���GQow�� ��S� �g���Ē�, m�aC\�"�j�6��~�I��n�4/^k[=\���N�܍���\o�ӄ�$ϕ����x�ɥ�S��X����fZ��U-����@�5(7�(~��� XO�B��0O���+�z�n�~�i$7����Ƹը�$�Z0p��]�N�@D���!5Y}��	DO�����!+}��� >�uq���>�l�]�/�~�����|e˫�H&���Eu��Rx ���1j��A��@���AӔ_�1G�?(��O%���
]�[XR�9�s,_U���WD�͘T�jڮ�l�c6�����{�����~�����y?��f��ѫJ�Ҹ�;Fy�6l���Xw�(3I�K�V����uuuup�����$��U��ڴ�Σ���)O�ۢ��O��?;?W�Y��>%7ߡR�c+��?P��޵#����W��mP��E�D����@�}\���`�K�$�����Hޒ���/5��/�~_�]8��&S��HExtY�L	�m��svsK���������5<kz��v)����ܺD�Ύ����÷��tqZZ� #ooĪz��U���Ve����bN���k�2��ڈ�M�I�_���$���*�ʀ[������ע�������e�o�Q��41��t�R�|p-L��nQ=q��jx��}7�@O3$���u�{o��t�=Z�>-9���ի��nh:�-՟N��������ʡ��-�O3��,��i��F����ꥉ���f�6�bX�\����R���w�\������*��
vn���.vO��y�~�E���n_��G����VCXZ�E�{�g�K���f����%d^"��<bhnZ��ī��giux)����"ݻ[�$K+��R\�������7[[�i��@誑vv�uz�|��5M��n��ɓ'�G�2%��enB���z��i@Y�;\S�#`�ߚ�(�m����S1���bc�fie�r_9�\ql\vl�AG��a���<O΋�g^�L�Ȉ���F��Dk�"�/6L�\�49�7R�4P
��aX�ee냂�l�/tϞ�+}��Oqk@��.��uf����D��G֮�g5�J������,�m�Qf:$&
H�6瑎{E��-��l�)�5 ��E
��9$�~AADH���1Þ�P�����V��
dbo�x��M锁����s�����'&�X�Mp�ߺ%oooG��š757뷠__�fД�CY�'?l�ml� ��ͭ���� A��z�*���������O���j����V�C�Su'��-��۩���V��e�	�S��s��'DhQ�݇�J��s{�[�a��^�bT�/9���WN�x���T�?M�ڨxנ�(3��8N���P(�}��B	w�-��+v�E'6��/fB��S�@�.�$��섴Od�V���$d��"x�$��b=]��O�vҪf�x�썊0R���J�V`���h�A�㘤�ۯqf���T�^0��;���:�v Ơ��q�tY��3HRހ���������ϾF�h ��(�������]�:5/�����V����>���n\?��y� ������}+M<�rݘ�v����ٯ���Ż���y��﵀m��}ُ�ŽC�nM:m�S
 ׮ن�p﹇u�ŕ�x����J3��s�,+�.�n�!ڏ�7g��o:�X�{^μ�vs#}2.������O�����SE�oe�#���ss`qO��Đ�q�z,�EşW&2]�L�\;�N_�ܟ"G7���$�i�8f�Q9=7�����L��k��Ҁ��o����U���VQ�+�	JLL4	�����u�*�pW@P���B#���N]g�H���Ĉ:������3u}���y���H����w�ii3-$�?��7����� ��l̽VPN[n��)>�"J�{ߴT'�q���V�y f��O�z�D]��<Jv�MOO�Q�F�j<� n�^���#�aD#	�p{�h�~h�JQK���_D1�4�����`�����;�y�+Sd��j��5�c>��WD���}u�T� �`��g�ד>A!p)�5��#���VY0�A���]7�ޔ�ێ�̭S� J��7Ls��u[p�N����i��b�a����S�w�!__߸Ӓ��ϕŴۮĜ�X��8;?#����� @��pE������Ju.��l�E*��O�)�����YHX�v��E�m��-�E�A�)s~^O���FCƽ�"o���YgZ"x����]�j0��7>�����r�ǏϬ�ff�����P�ɭ-��t�0yD������X)�%��T�Ǒ��b��2V�t��l�X�0]W���Q���=A�O-��q �\h&�[�F��Q���G����,q1��hx�8�/9��0Q�K,}���FE �)��ޝ�#��8Z@�$��S��](;#0�E27�ۗb�EbK��54BΉY� �q��yx�޵©Y�%8���c�gc:"4��$	��%�w~��X��sa1	{,���N�ϡ����'�ꊋ��'q��Pwl�!X-��5�Gv��A?�<,�#g�
�K��1��hos��UM�ۄ\y�uqJD[u��9����+�Jb�/�E��0�� �	�˒����|6�4��Hݙp=1�>칯��]���'S0�4Y>>h&��Q��J�HH^*���t�M��ߟ���Qw�Ο�R�a�<��f[0ؓ����O��c'�im���5P����0|9�*�u+��ND>�s>s�v���pB��W�f��)������X	S�|	����r��}M]�L��w�>���R,O��>�˝6��������R�����F�d�����^k�*S�F�W�{��wddv�i���������;$)���������k�N�W��3(o��Z��<������cRYx�U�m=�x��+℔��襤e;Z��>�1_*)��n�2R���ݖV�����*U5�gnm��)�G3@X���]g}��b�>�M�a��%b_��ϥ�!�t�m��<��:��?�|����p`�b����
[X�/*�1,�x������/��ܲ`��b�{��;�P�׈�Fp6͈���Pw3���G�s�N����?&��LQ����v3��D$e�w��FDI�,�oLV��;��:P�}�8b��4>9ە�f��JbT�5s�v�B����ɂ���]Dw�����w.7֎�յ��\s&U|��l!��n�:�[��I�9�ŏ��ʌ��3���d� ��Jk`G�U��V'���pp!�o&�^�Ǔ@���Fb[��&/�1� ��][�� :�ք�]�\9�V��5�����t��w�\�6詔��,Hs}������p*s<!�:�\ܗ����������F��灭.�<HG
��jq���$h?����v୬�h�����R����u�c�
���-�&�,7BzS��<<S5��/=��h���%�'�޼+"i`���0��z.�!���N�ޱS<��m�B��~����Z"�pe$dI��6����۾a�Ԡ��+��S�5��E��OJԋ��Y��I�ܔ���V�@��'�0类�c��G���ʠ�'^���oV�,Q��E���'0���a��,Z��+li�X;}�9d;A�~���+�|.�w�� Si�譀����ޛp[~P���Bp�n����`i�$G��{N\���|Q�9A,	c���)����٨x��f����V��M����I9�ſ��h-�ҝo�f��k[Ѵ�����7�Eb5N��Ic҅W�	5�n7ɮ��9�j�h�C�ަ�')RvM"J9 U~�hf�z�-�g���K�+�}x@j��L��J�v(�|� z�8���H`�r5+��>�J7�R�����!��H_�-�}~q�İ�':��-Iv0_�L�_y��]��r�{I����xtd9S ]��\C!�_~����V<���T��r���Ы����R�=(��zMO���qod{���"���8\��U��&��p;d=7	��I0T����%3�[LK�8�I�<e��lLkM�ޏ��������R5]$Q/�������e��%1�f �nz���He�� d�u��գ����z�	P C�9�a�yJ��ѵג�%�=�w�&���^��.���_��@�l?Dq^���\NbL�z������p���Q�<�[����_L�AGWw�t�oeu�AL� �9�K���M��{L(��-�崉��9����k�}Px�{�;t9�i�����'�����M�7�+P +l�/��P>8U&��y�#J��h�ݞ?CQo�I>���9d֗��3�8�	Vf�w�[�3�g���K��tw{��p�`������\�-s-�w�@��R��v{����x�Ā���Z�`?�y/��s1cڿm����ϖ�H���MB�,�\0i)�ۘSP��D)�~Uզ�^h���dk#��^�^�ɼ۹Um������	~����i�����ȍ����ߦ���)���͊o3o1\o5M�ر�m��kMMu����xV�����ߍkކ�<]v��N��ѻmwӡ�1ô����}G؜��m!B���	b��Z��OC䢢���@�w�P�s1�mpd�����HC ��6+q��e��M�����"LY4i*��}�����{��Xt�U�n�yj�HO�#̋`���M�	�5�%*ghNO�]%ӠOW#��\����]ڡ�0��7J	���X��w>% ��8��: $D��F4@��!ig;����E]d�����7�`���+3�Md}���2�
|<,�T7�U�ҝ�3�9��+^_?
7�o��-��m�I�)�C�8�MqA�.���7L��AC�>��W����tʳ��me�[���=4�?���^�(:�뻋����ղ���2zJh�p�L�nˌ��=�p�Y�tϕ�n�=p�����g/o�W�g(����y�zn)�j��j��:=.
n���&�$��n[�K���[_���; HwJ� -���!���%�HH7
Hww�tw�4Cs�������.�Y�N�����>����_��*�Zߚ`�PX�(YA����"���a6�;�&�����!����(lޏ��5�����N�sۣ��e }оOB5��&hk!�kq�~Ҵ�(x������918dPu���g�:�V���Y5�3B<
mB�Z�� k�/h����8����
@�hN��t���&H��Y�?i[1I�Qo���ov<��_��B?�
��(n��!9��/gd�D����3DaSr���K2R��-�
�F�A���sR:�M���'+�k��s,�W2�~~y�V���Z�ٸ��u�N�%�|-�?��am����i�����v��m0��"��3��M�P�R��M3X+W2��VR�	k�	+��'��\+������J��&�ļj�x:��� �i�+'����q�8��R�J��.jh\��v(�s��/�E\�pE�,�W��e5�P.�
�SN��T0��W#�ʏt�E�yc
�5C�X]��S��	�����+.!a����QT^..#��;D霒������Oi7��TT�{���RՆ7^�zEpq����i{  �����Sa8,R�t�ϼ�3Ƣ�5ȁ��L����+;?�%ɾ�\ZB-4:R�Q�~�� �Z��ͼ�ԁ��!����:7S�m\\7���a0Z�1��A��]	���;m�q;̮fiV��f^��W8�mO/��W����!�"��A蔥����n`� �ixV�V�X�fFh�Z�ͼ�{Y٫n3p���DO򪨊Y[�L���"�"��@�l)����U�|++���|�Vpo N�H@@��N�ΛqI�N �N��� �`�j�&����#���	 �-=P�ðֆڕ��݉�%�o�����w�j��iC�tCL��B���Pâ�P�Ն���xXl��Xɀj�*e�'H�` on�P�����3Q8ɸ�U��T���QD/$���h���w�c0�]�=P�9h�q8YC���trv�.ø�V�{Ҕ�`V���:��Xs����4���h����&&�,+ˬ�a�����Mƈ�tk��r�ۑEh�\����GC�̢p(����6�$h�U[7��j���n�>�Bf�yWm�:ʀ%)YO�����շ4v�ޑu/)>D�-��S/��xG��)~�?���3\�j���_����F��TU���&o�^n��:_�҈)m�4��J&MK�M8 �������-�rc�
��brw��A�GY��؅8��&/�穰CRH�LE��U��?U��<��|�������aJFrk!��v�<R*~h�
]�ߴq1\��e�]���io�ʯ���iQ�s�����hʐ�%Xf�JH�m����)�:��9
�W�?�_�nʴ�����C�{�ga �5��^��ű����@���ox� \���� ����r������?2�`5-����w�a�]
[q��{u;���,��r�����i�F&��='n�q=Ao@��'�����w��r�*�F֫���o|R����_�1Q�]:��eaŶ@U��q����TV�qZm^c���YDr)ľ��P8ު���o���o����"w����R�	�]����W!�7���7���Z_o�Em����6�^�C����m>��
�����UT<*����k�d_��
	���TO���|c��yN���BW���R_���K�%�W<?L��[�Efe��y�X� ��p�x0��JT$l���E���V�����2��|�s��3�#�x �]ޱ��ˆ�˕�>�����*���*D��Nl�?�u��s���0N�U�ِ_�1�
KH�1L+�3�N;;S���;5���M�B��PK��r���ά��W�ћ~�ll��cjJ=W��T8�:�A�
�»�q���}��"6��i#
����JEny3�pZ��4+:2J�e Y��ߵ��N��A�!T�J«�#�z~b���xȣUrr�3nfb�����b��~�5��F���!O^	uu�rݖPA2I*h�yr�6�gsP���E�4�*����0�A��8��g���o#M$h��2/��thZi�Rx�;|��f�
*j}��nlR����
���-ll `�/}�V����F�'���Fٔ��_+m��yW���E�P�*�>|tx7;�/ /�k)���3�z�+��~̳���5����`k@@�<��෗�.m�p�{n��.�t&�֔8�y��mG� ��ő������xdҬ�¦�������:~��*O1g]���k,΅ҁ���
��jL��q���;\[�;�,Ns�^ۿ܌�x�	I���߱��i�嵥>1' R��ѕ�%'@�4�c���Q.7*G^C���yqi)�+����j����(��+  v�RQ����<��H�>_6޷�ɛ�^�^�§������9>^�Y���b %�J�BFC��t�<�$�����-އ��`����к��%In��a�V�C�k�Mʠ[���0�Pk����<���P8��Y6��h������hT�hQ�ߛ���Ń�����հN�/��9]f"%వrLۗ��;�8�E++��u	���j���=�R�]��Q�>N�e��7�T���E.܎��BH���[���v�®�����Q�@�Q�連�����m9�ߕ ݷ��z��`�\��xSu�r�4ajV�A�Ѭ��O�k;���w�,��؇������!��f�m���b��P~�91��'�Ʌ�9�B���� �;X*�d�Gyw�ͥZ�e���;��8��)i�����=��QCh&��<|��҅�R��B������yc�#��}��)�|�_��-���H9.(�D�16�>�������e@���59�;E�W�?=WK��F«�g��dߡ�.����@���J%\��54P&J綴�f��8"�I�]�T�<(`���	���n~A��9S�<�,�QWW��3^���s����~5n�i��y&���s}e9��f����H�[��(�f��j鉶����zK��64��s��Q�)W�����=N�1����gϨ|`onXsI��ڹx�7Vie'�$�.Nzc�V���q���Z�3�ۑ@ X��.���ר�¡����l�� �5�������:�P��t�t<�(�et$�����^����j�}�qqIH
�\�2�'O�f�GI������2��u�n�SPЁ���ZRn��,>AmBhn*�Y_��Ѓi>j��Utd]��D�a��X�'�d�gw�s؇��F?�Ӟi�TE��q[��f�:��h��Z���q'�&�� �=X��Ք�," �$�vԞ��{�X���)���=̤E��, پJ�����nj�V��������c��1�^�A�3=��{��X��W((��s���Y{��?4K�C78; ��f��LUkF""�y�.Ӫ+>�_[9oi�	CQQS509g�֌R��o�=����K3���	�̛��%!Aѥ��O<:�R����_X|A��`�Z�a�+�Ģ��3�|�II����4��m�F�9 SPP`�\��4�)^�x�J�_�>�[gX�U��uj~���,I�_Q���Ph���}��9��k��AM&���7���x��>M��f���C���gm�y�.f~7�-VE��p�F�Dѕ��������/�N�*((�������) �����qXwC{������w6��G[3����JN���	d!
��,�Vq�o�y~�x�P�0l8�g�d��F�.-�����,���&'�8�3�#�bJ�-�"xYy�{�Ru��y���@b��.�����b�gp+Op��a[��m���W��X[Z�s2��Ni&��6�!�7	VW�� ��F��$����7���մ�w@p�{�t�7�ao�?���C}��j�V��Q�����Gpb��>�{FvտCdp~TDD)�ϧ-<rUU�'�\�B⏸Xgf��)))7
Q*�OI�q��,�@,w� ;d2���>�` �@���n�Nq;Sb���p�91`���?�����/@4�{�l�AIJ����ͤ�#����Z����4��4l��|^��n�,�7gy��M��LL(b|�%O��~��<�a�<���$M[��F���~�.�L?�O_t�a-���~:o �P��h>� �+u?X�����(�r�w�w����tE���A�rrr����ⶶ�¹�$h�2�S1��:דV �e��6��e�Q�+�f�~v_lԜ�k��4'3o_Ͼ�O@Cvwߞ�ޚ��H5�o�Ŷ|!�}�Q,*|/^5�|��"B*<n�[Nb<�rCΥ�fF�x�=���>�R��Yo~>���Y S�+w�|�0~lY�U�`Z Ġ���~zz�M����iH/�z�c���p�]�k�P����#m��{��pbd�l���D�=�J�$HBR}��_P�1�LS�=���0J[G�!�
���$\HLV{;�oiqq7�(2
JnE��(~p����������{i�m����#�@�%A�?)��>X�rs]��4 �w;{�{�|�,��b���)��tRxZݿ4<_�������i���Q�5�`;�J
���)�B��暸�`��t��!����>==�&,�F]�3�%p�d�\�w���J[��탻
^��F��i�k�zLr�U�y�.�*����=�j���B��Z�"���Àn[qX����ov@4�A���^^Ҟ���#�+«S;��;��7�=��(�d�:R��76�hi�X� �_� ����- ��9F�.�t̩��3"�ĵ�x�;S@��:�X]���Ӡ����04݁Kє�Ax��Iv�QG���`P�XT�^�s�oP�,E��@�x�Cl�]�����.L��8�~�1��E�da�{Ţ	��2]�Mۀ����.����-�'��۫vc�u،�g�/Q:�6~#�J�ZRV�6[s��]|9�>�i+W���NN��`^���
�@����7Fff^}�_�;1�\"��O�<j���/)���?V�-�o��b
�����>��fY�����C�"�/�v�s���Y�Ч���k���ss�}q=[|Ŏ�7�K��0	��o&��Qd$@�D4�� ٓ��!��瑬���� ����\Nm]W��C`�h7�v�d�5�pm�v�'ztt��%Nؓ|��6Y���4�ȩ�8�?߶�=PJ�ϱ1���Ϧ畒�˲_���,l�����K�'��ɚ�k�:-��rd�`##�f�ss�<ر�P�ORKv��fh���N	�>���y�#�F�[F��}���G*����r_MW���Q	{���=��׻_B�����}d�k(9D+'J�`^UU9�_[O�`������9�A��@Z�n�AB�~ҫ˷[�A�#�;�|0��{�0H�sn�QSe��gf�`�A�ӁT�~���=��i6�H�����k�¥DFQ���l��y����T8��T�A�)�K�c �06������@L�.���3�����V�Z�y��>��E,��{�j�}�.����@��q\����E(�:z�h�M�&�ȹ95�6�,s�}@{�3=%]٬��S'H-��
���$Չ�
�s��:�O�z����ܭ������;t{Q����$�?M7prr�$�*�b�v%����2ޗ�t.��@j����֊(�L�'"�!��t���������;�]���m��p��zG�%

�큄LV�+�,Y����bO��'�|s�0���7 ��d@J2540��c\����( �6$>��p���)��@�>�-�O��O:�?o1��2�D�5W��(9�o�"U�[������㫡[Mnl@�_ʽ�ȋk��)�2��s�1� �w�du�$�"��I��k��%���D���ET;^�[ߎaPBs�f�=������V��Ս���.(Th=�;�.�6�{۞z����VV�����0$�1]�П"&��R���@����ȸ�'m�:D��z��Q��(QH1��mB�k:`���Z��u���"4+N���|��M!xz���۾�W�s��"��W�e���!8$)��O�_�J���!���h�:4����n{�ԕ�� ��[�x�����=iگ�s�9���FQK�����ۑ�Ԫ(EH����ܩ�u��i�x�F���'�Ԅ�~9o��^)P�Ȏ�}�@fq�0 ���w����1�&�n��M�L�Wn9���+C>��������R�׳/G~���١��X�~���
n>��YW� ����imܭ�������6�� ������2�%�]MvC#���=�Y���
�HW�����^��@߿Wf�)��֮[$n7
�'i�����D;KK�$�bCT��Gd���uw�ە�'�vKz�ː�Ușk�r-�O{;t^�Tmwrh���Ki6cY|H���#�`M�%�oS
zX��8�?�hh�Wy}�'�@�8g�h3�%H��������8}bU��clr�yJ\fT9���5�hY���MSH`�U��p=��d�q��ސy��&V�
b)� Æd��t�|����mGPg�|��n�psE��8Q,��?gl%��z�Cp�Rq����dB1~hV 屙�ʖ畤���z����:�|���h�-F!'�d���IB@02�K�yZ���3w�9��Dk�cخ����f��`�]I���Y?��c�b��3������Z�yO7����Y��������'�H,���"Ʌ� �W[v�i2�(p$й��=���~�G-Aɲ�XC&��
�b""|ZZif�ʈ�;;�R�2�i����ǽR��ӌ�\�d�6���$�+��aP <&W
��6��z��'�F���Ǫ`)���T�M1�Ց�ÄG��{�dai@k��2X�\1�����h�l�j� �^u�4
Y�瑟�5qY0>���?�H�&���>@C�B��@�� �S�k�b?Ӓ�Iߍ���G��lu�R�kB�cIR̩]�{��r�hM鼞�ϊ����vJ��"r�]��>ce%�K2��A!���4���QUͥ�^�f�fx�G���P�`qf!⪪J�>Պ�#�e�i��<�h���p��Y�z�m�����gTl��h{墙=i���ϡ*Ŝ�]���#�:m���0�]�EW9+b����D�!�����{2��
Pd^m�7:�e��Z�ړKK���ϥ�='�s�_<x�O�tZ'".:!����
1�h���]�Rq��a�]z5��S��m�
�0��%�K���!��ׯ
�G�_��8ٷP����O����E��Zb��v�����M{��V�ᣧM%��L0r��o��țy���1�[��\X�T�II�m7p�S��F���j��v?��&����7�F���K�(��5f�l�j��͉��K��ȝ]F����W�f�GV&�F�����=Ti�Ο���l�ina!^XLf`�8c��ta�q*_`K��pg
�y�i� �	_�6�A�*z�ڥ5Գ�����;�Xc##�PC�C�@���*������'�$�R���z5��.G��6�/(�J����E#��D8u��X���[7���;wO��v�����t@C��WR"i����CG��$�Q�@C{�"�)���0��܆�l�"�;��g�n�,i~7����z��j�����P����\���ۢ���,���m��a͢�;�Sq+<4�$�M~$��o�)sm�O��7�-
j��~h�j6}��x��>Mկ\�ؿR!�*�d�J�{��� ȠZD���hf-�ۧ�V6fD�
�]�ra�PzAD\�RF���.�?������k@~N�C���B��5�IvN���������9H������H����6��k8���7�֛qr�������L5���6�.����~�r�Qy�f��U���:�eo���.�Gl�r��y����KhTF��%>��{&6�F� <@��͓#���w�����C�t���q)#�΂�����B�L�7���?|Yc}U���Ak����"�^;M���ת���~]uޜZ�3b��)��1ټ1Ċj�*�wf���\���В��J��2�je:�I�\�:r�b��=ʛB��h���]�c\���2$3MqX�������f��|<��˳������15�9$<�t�ɥ��B�%���9��
M�gp��f��S�ju�OS����w�f����?[A�?��ϔ��b\Y�=Nx%h�<�+q���MEU��q݇lv&8q:�W	%���kOz��;.^�Ŵ�`�wHE�v-0bY~G�%հ�pA-����6�z{R�aB�X��@�JPT�y�a*��h_��\��6�f�K!�ES'����ukM(�\%�O<�7�^�.�l�������9xϓ��Z�������Cf�Ǻ��+@i�8FG`W�*�/~B��o�F|�=��Cʃi)|�0Z;���@ɏ4����mV����ɣUn�3��ϛ�(�C���\���sq� �k��רJ�C�.�e�_3h�.l�$t`; x�u���t������?L�_MW�/���M>R��
��fl�|�X����&��s����Oa,�q�qQ)��iW�k�d���f`al��Y���ipWP�f��4^��������[��{$�B���#yx��`��� ��b���7I���S�z�z~O�Q�ц66G����p�A]���ذ�i�JitR�l�y7�������-7�5��˓��d�Ͽ�Y.zH!{����ӟ��qOv�* ����l�� Nc�o$jr/$�+�R��iC틗LM��ǎ7���a1(�c�N-	˔��j���@����tT�)�糳��7����-��j�0\���33?o<] �@�w�m�}�fv9wwpk��s��QhL�OY�{E�+K��&�ї��Jۥ�_
���o{k�'�oP�����<��	A

��{�n«x�)=�1�/�8�Hx9�=KU]l*�H��QX�jg�L�Z?����;<<T��T*w,o�,0���a`b���O� z��kr1�P9�˪��b��7*����cE�����EoNGTT`��8�����M��i�@R���e�B���_�a�K�Ԏ�R�����D����|>�Y0�������F�_��B���gGF?p,rv4��9��*�/"���z��8��oq+��5��\��|N���LRpEU3�~��5ʗ��_!�nza��( s�*$�^A�_�+�n�T:���~E���Z�Z�	�<���]IT�c�i����ؚI��>�4��&�ƤOm��O��M�����B�C��Iy9��nZ���r�>�??�����o-�lY^�P�-�ǜ����tw;�,]�b`<���(�3-u4��~y�G
��/�0)?��n��J���,��'�R©=٬�y�/E��?�d��X��ç���UqN���jI[�b@��9娇���SڱhS�#���N�$r����?=����[��/��t+&AT�|pt݌�S���+,�xD��S϶�?88b3Z��)ӽG7� U���t�q�f58�~#�0~L�$ǌ��f̯�I�1
���G3�}�,�����]a."&W�i6v�D�_�X.Zn�ý����6t����J���%�&Pu��E���3䊸�x�ﮊ�G��z	�G%�,�u���M/)a#-���(��Kب|���2c��7�U���{��@���_IB�0J�u#}�'�G��H�����xa��(2��=��^ZZTݗU;fW�o�$#���'��W?D7s�l<T+��@�F8��Kr�4C�!jhL���c��c����cZ���F\*��DL_��V�HJ����&����v�Q�+�iO�熋ھ�(�+��L��h1�sm�87�f*�qeӑժ�Q����T�R�X�>�	j��dZ����ޤ�%Jc�@�}ۤ(E��&.=��oj���¥�vk��n ��G-]^0��{ָ����S����.T��&��x�0r`�hؔ%���z�K�(-��A�Ż\x����-�������$��L�Lo�{Y�x����Nt_�!�xd�� t@ŇS��9�A�L@�O!� 7��!`A�ݎ��vlXI����cN�nV����)���E�ZU��H�ɇ/�����,cU�θ��OxC�v�F���/��÷m�W�`�p�Vp6��L-t*=5�p��Ƀ5��=�����$�:ӝ��j�"������P���/��JGK�ʥ�ӼMc���6�ã*q	�뺊͵:�9c�Ӧ�*�φc��������L#,��M+��_�ۻ�[bH<���E�ZхG�9;�׼��՞$����>���o�\��7��|�	�mm��by���K#2L0�Cc?��ӏ}���a��%xv��u�x����x��i�C�uɦJ�� 2**�;�(U�jx���0�݌v=�B�e9���E$=ts��u;��vIK�����+-%�1zɽ�Y\0��~��������W;�u���g]��3
{Q�����6�
�B8��I��%��4��)>���-�i�V���BԴev
���3�_�(Ȫz��1�+���`��0z�{7�o�f�fܽ���l��+�9�)�'����0^��}wH����
N}��y�=��mB�7=aJApVM�x�0�p�Ĕk1��m��>�æ�����a����AN'z���P�r��?g?��jv�o��Ҭ���X#�K�A�Y�E���zjq�i�/5��h�9���(�'������Qr���Ip��=�����U�k+�	k�Z�H�T��ɑ�
�oB@c�3,+�.1|eb�0��o�ϡ����OMf�ۡ���J�園0tv��i2��;�UM{��>V8��#QB���t^�j4����*�:�{:�wxh��Č�bs�
-�qU��%�hs��N��$]��h�p�����,pN��e�[~IDm��q��`EU�m�,.�ZY���pr7#$ 0r�)�1^������=�a%c�F!�w�d����\�괲ξ�ǳ�#��z�[��+�\tʗ��O����ߑ����w�F�X�~�'�2S48=��&��Zh=�@I3f�h_�S����>H����y,obs@�y��t���iM}� �?(3�zxt������R�M�����m�s�mq�"˓�׬X>n)`�uy_�ά���>�C{�3�+6	#����^�v�WP�j����ά鍕K�:2ul��@(�s��7́�����,G6�Xx÷[o䡰G�Q\V��<&ؓ�݀!�L)�ruu]��S-�����LxC��.r8$Av�k�p��P�����p���H��kǽ��2�<IT�KU��n�-mJh k��g8�R�w�rt�A\9�)�h�˱��ԥ����<��2	�^M�!Or�y�0Lw�z����K�!���d#󬗀��ƾpo�#B�k�b��}���X���>l�w(K=w0��Fz;���KT�������>���|�.�M�+'wU6�h;���j귙M���� Ł<�Բ[%��ԋ��EIF|�S)�;U�s|:;e���nn�"�`��b����;{1ݲD�w�zb"I�	t"r��|<�:���{�y�r�c����\�u��о�br���r��qv�������D)��� ?DP��s��d�<©	<:L>a3�8B�*M�|����u"'B$$L6��ܠ���g���qɎ�%J��dW�Q���*��<���V��3A�D�R�59	Y8e�뽧.W�e��(z�}�>,7(;�Wo�`��I�]�}0罧�� �\ۡ�e��l��o�'�E��E��:�3��<K(�������л�\��%䠝��q�R��A�r/^�w�K;:1%VBbLjiO`�4f�ƣ߿�;��wS.NX���l�?rQabI�Z�f�y��k�w�vHZ��Ãcy��:���˷*�G��7F����g�y�rY�Rv�c�x�DO��.�M��W�Xh|*����_�Y�7;\ӊѯ,��"�������b����]2Lؐ�#�-~��*GO"���8�H���>��h��C�<d�5Ӂ�����<�b�<���<��Y��Q{�f��"����U/��}&U��뢓.�.JJʃ4��vm_0X|�42
�j��aR�&`�G"�r'J�P�Eva�v	5ɘ��e���(�Db���b�l�{�BCy���~����,�X��zaKcd5��kY�[<��k'�ѩUt��o�7ihU�}?D��p�ȁ6Y(�L߷骪��q�Z�1��lIyyy��Z������c!�Fjo���98���@O+��T��^f6_vO���}�c��95<�ˡz������v=f� ��uM�����yE}cb��d��&��(�'��WZ�l
�<�QQ'h��G���*������Qb�[�-�ji�O��7P?>�?����+�}��RQ�;��pkA"x���lqq��R�:���,�|�ivU��3p���G���g7���ߊޝ�?���� ����ɴY�N��l�����H�-�u���2Ɇr25GTok��;d��c��P�~f��4Zi�!7!F��U���#;6��_�C&0�c�W��i?��g���$��x���V���IV��Gxd	"}$+:=�ĩ�6�vq�4�U�'�'��#77��z.g�q��#�<�y�^NF���\Y�Pg^��zί�#�ce����~��4��nn6�}��8!�� yߧ?��%�+X� ��f���82���]BF�v�۫��6ZϹ�)��M��.�o��<�h>�������� ]G^��6���ه�M�.�R�Q������k�[��m66Q`�*K�1%[�_��3�p�E��,�ƥA7�k�F�t��`6'}A,��^y��j�5�>�����rk�����])�έ�Ǎ���������=F�!t�l�?�d��X_'���Q�O�4p𯵒˖Z���0C,���(����i�&�U��c�5o��0ܕ�O�`�ȿώd1bL��v5r�+�Y�����NRB�{�z��A\0;m.�o�s#D��F�Ï9K�,����azn����'�� �B�V]�<f'��m]p��E���������=���+� ��I�l��~�?�k}լ�� �V�U� 'K��ed��Q���x�JlD����ddd���h����c,Ӧ)w�~|zC*��U������S����_��c�\��J���a;^.>�չ���t��m�y�����lS��r����SApϢ4	��#��{�7Y��^������I�J$�����u��0�(�"E�Ꚅ�X��s�M��E�d���_��\�ݝw1^���)�$�ώ5`�2>i.�mb7mZi9-��z���at���q��(�B�����ϑ�E�|�ޖ�s?�=��qa]_E@��s�b䶵��f�1.4�u	�4/�~��6�������Cӱ�$�
9Gv�=�*�|Ś
�}�
�E�����J%݈��.��	/},S���lvu�0��/8I�F��������O�/>sY��� 6��vue�� �qVچ--pح8����	�o	���7��lQ|���q$�%A{�9I�$�]v4a��K���+.�|�z��<���~B��ƅk�����&�f6�`��תt-�EhJ�1����w�
X`��x�� �ؼ�\ ����{�zV |��7ˏ*�g&�Ĕ�ᠹ�����_�d?E���ΰ�.���Dɾ���˩4��JKO��9
�lRecK���Rr�%���C���,����*��[��wdSJİ��v߻ZKe��<ڿW���X����x H�m�HH�k��B��A����lr�ss�x�0���H�)�G���L&��jW�S#{�X��c�@C�B"�g@��r�8c�r]�{YK��=B�:6
Ѡ7����2�-���u[<n�ߐ���fq���hPz�,��I�X1C_�����V:;;K;�QPQ?��Y��(7g"S6��D��}�+ۓ/�3����S�O��fw`���7M9G�,��T�o5�~!�8�%���վ��c�1V�&g>]彞Q�5zs�س��sh/�^��{��h[�ޙ�NJ���u�K�M�HY��	ЮM�L9����}�F��&�zgQE'���~ܡ�F����֪]�)��Q�d�F�}s���ߩajXi=ϔ�{o	*_�OL������2.��w�1��z��:���3 �1�R�$-����X{]���~ٌ����W^	[����e��,Uw�-���	O.����{����~�Nt�n��GtxH�< ���ؽ��~O�F�j��mo�e�ᬀ�G�s�ȨF�Ҫ�����0�p{�ē\��6|�u���Ғ���|%�+ސ͘���-V��:L<<<I�֗�f��_���9^j
2��G���I 3�����Z���Ye��̏xg�b�YI_L5a���P�m�K�\٢����>w<�[�)��PA���<T'ڭ��i#��s��H�u<R�^[�Ħ�U�8�s/��ڏ��q�7hh�3�L}��v�iΊ�����(����� ���[ب�Tr�Ĩoj�l��5����=�/� �6uc�`��������W�;.���X�S����F������w逘߽r(����E����8�����FiY���X�!�Ư�u���'�����j}�����BB�$ �v;bL`z��~��UUS��C+O�Vp�d��
�o�=o�}�nJ����I����z���j��Yn��{/���1[�&K:n0����k�O����r��~���KF��Nq1Q4�?�8!�'|��+�:�b�Ue@�<���^���ǽ�$��'$���^e�{pm�9w��M��g6�� 2j`q���$z �=�R��0U����S�ڛ_q�NM��ur�\%�ZJ��5����ep9�ޜ����T��0'EUUՉ��cP ���x������7)(�tgd���O�}h.�$��`x�@�c6�·��7�	������vL�B�544lQ'ҭ�Y%���ԙZ=�77����h�F�M�� ��2J��w���&��Y^Nn�t�"�c��0�c��W�?t��Ca]{���.DX�cX����T���.5�'���8��AE5󢷾����7J��+��*���G+�:����~`�\��d���-�yf$�^��,)�^ir��p�X�W���o0-��`YN��ׁH �@=��:��[�[�{���(��	}nX���xXSW�w��l>�����9���PU=�������nbBq�\?։�>6,L	��k��֖�;%���Գ\h�,�F� �?B��g���2�7�bh:M�-��!�I~!^�8�O�E�ܸ�CR�&GOUuii�Ң����ۋ-x},�Y\B ��#D"哦��:+���O�|\�؆��C��[|�?�P�8~6����\d���=>p088�V.�&׳}�-^TR�����2畆�t3ı�Vv����A\�q�,ȁ]b6`:��2�w]ͮ�I��v����B^����&ڂ���:���x������"��Ӛ>L�ڦxm�қ�t���|��rW���~��j�l'YR��#�Nr	n'�������Q��:�j���9�OI�	y��=8�����2���������Mzu���	�
��/`}���$�Pot����)�[#5b����ﾼ����K������b�8�J��)����n��}�f���F�Q�tۍ$�L����:�vI�d�0+P��O�~11F�1��h5��~�����/Yث��$"++��8��G+D�{�+��Pg�����F/��fgX��I��I�/�.����@�����#�5�~,6�h{7�T��=MB�/�� ��Ll����O�x@��_�k��&o	v�[S��ڻSS�+?�
(o���˹��k�� E����yY��C&�^ON�μW�?M[�QN�9棍4�E:�������?������&�����>�^j��W[�R�/�Z�8���v�r�������\ZN �����$���4�X!��"��v�ہ�Z����N���h%�qd�2&8d�gh�U�?��/%(b��/�09XٴVغ�w�~��U���n��
z�-�I�Z�-����0�ޕ���+�������囿�3�q�l�!/g�]���_�?�2��I=��c�{�ʹ��`��_r��!��gp)��87{�XؿLl�v2��t+K�/**�(R�B��2��]A��Ց1����iSG�|$咩~�ː����� 5L�a�ˉy�������O.�.ʓ((O���[����k�WM!N0.bJj.,˿|�O��|
-�������%Z5��]�s�3�5��n���-������טp�K�}�3�~ON��)T����^�YN�|K;ѣ��07���7
%� �w�$��m�$P��8)�2:���$��� �/�vyʇ[�z��++��	�V�Je�ױ�䥟o���k��©Q\�6;���W�"�]c@HM�+׻v�Ԟ����|����*�ܺ|�_M2դ��\lҼ���vé!�gZy3���?t���xs����M̠.���L!=+�͗�}��A��:����aFiU��bS_��z
��A��oB����J7CI_RVUU��~�M�J�U�ѭ'�(���M�ΪN����~MO#�3M�u[3Ʈ!���}y�)������@=��3�3��p氿��s��<����w��y̷���¬��"Y��5V$��&�X�T��[��#.@���^�&��I�����}/���:�=�ݘG�����T^�v*)�܋��ǣ��{�8,������������Q@Z�D@�;������{)Q@@@D@�k)�na���wQߟ�����sfΜ�<眙1͑����+`�-ѭw��d��'�7[r��g¡abn$~x����9X�I-����r�/���0����E���$��P�͵C.�!܋�H_�VB`�P�}�Ã`���kH}��@���u�w���j^P��&!`֡��^�2�[���7�aJ�Z�UG)�gdg�v�Tc����S���X�g;+��L���/(�%���Ř�+<H`�`&	=�����lN9I�D:m���Ϲ9H���e�`;�,�($��L���xq"Nub+��J8�Ӹ��f�ax!c�)n��_е���C=#�+� zY~�eo����A�IX�]���a�B�]�ow����D4N=��Q
���6�ԛ�������$3+n�T�/2��� [x����F�*#���k��[�6Q�sx�=Ӣ�a��i<���|��_�������( *��&��W�;��NOO3�m �b�e��/�����w�gc��$$Jw����S�ѣ��A�'���"���E�F+�WD�o���=O\	t*צ�ʬӅ�T;�cdtmA��F0O$�rJz/S� ����n��Tf�����ӭ�1`�����U\�ňX���~���\�v����<U<sx�,\'��
R��P�Ȗ&��g�@iw�%jl:f�a�i��i\d��.��ގ �
FaƮ^L=\y8U���-ҿ��z|�������Љ(���*��;�;@�����y|��OW�<c��������=Bez�a�緑���<��ѧ��en{3�ۖ�AAA�M��[�[����W��r�	��;7-t��J8��"B���TfdOC�k����aFu�uq�"~c���i�h�aPќ�_1�Mr5Sf��pKq�5Bbk���0r���]��EoD�UA0>ρ��1���Ի�.`?ջ�B9���(�9F�>ey��>_���ֽ��3��.&�NZ��}�!��F0�������;�覠����#="�^�x�e���\}�G��yus�P���0Z&��>���Ưn"�F���$>1]]��g�!M?�wS'''�Qc?�lsԁ9�߹�!Qw�C�l�xl�|��t�D8"Azh��&���Pq
s^�����0q\|�]�*���"g��TB���p2I�����ל� p�ue�[�wE`�ˁp�M�%�U��a�)MK���X�
�!��S���>,f�H�{0���f��a����m��҇�W�"��o�h�(�5���/u���0���b�M:)m7�~�-<@�^Ap�[��*�iW�΋� {/��a��}���3��15�9u��V�i�R��e65!��[�W��}���+���h����̓�����v��.S|`���z߂�4W���'�8^b��3�w���$�5;��'M�	�@�6�$(hh{���|��54|PDq�V$�(Ace��K�Z�d$���J�&���L
P{�fc(���,_	��i��>{
�Fm����.c�nP�BG��Ɓ4�V�����F��<l��6l�S��4V�)��k$z��{�A�-�[����Z�#�cJҧ�������{T��-�����ߕ>7%���6�����/g&�p�dI�D{��gk�����ئyV^�'�_�9����b�v�7�	p���E�
�~K��G��2Í4\�耬7�S�����n���]���>ל>q���82��L�9�u$q���\�߼��R�,F��Ȋ���R�vω�-+�DOȱ/�Ħ�3B�;;�yP_`��Z�,��2Bl����G :R0�"�%��v���4Wi��Iw��6��p�{�5�#"\l#sw8�9hwnG�#��Vɕ"n0��&�R�`!���+��.��8B�n[���k�`'@�TT>�L�}n'��!OF��׸Ε:%�&-sU#����_Kw�ߋQ��J6^^)�h��b��0�n������kT����Rވ�Sۗe�e�k����bj7�Ժ'�����S���R��:&��ƋJ�h�$߱��mά;P��FaѠcf�?���y�����5ߨ���{�9���
5g�39XxS���]&д'�Z{���ʘ�`L����Gj!��{n* Й��ӑt��>23Ӗ�U�3S��b�G��\{�n���^E�rK$͒����kD�q��/�o���\�rN�S�[�{�����Ƴq�����\|]��=����t$
��L���?��p{���c��/d�(dH���lstei���cv~^��ϟNN�ũ>B 5:̂�)/̐��pÛ�|ۖX�m2n���l�-�U�9G�yM��;]��S��������>֭L7xr����Q�{4�ͨ�C(Z�i���ĒxT韵�t���	�i�����:�����_�%�o����i�gr�2�	��K�>�C+yO0X`oo������p)���%��
'�s���0X͆d�g�a�L1R���x.�fS���nu��_��R�5b;Bph7wv�{c� |���AGg�c���΂��;����>'���@�ۤ�e�Lg�o/-?~�hbU���Fu4O�Vx��/���]F3��� T翠��7���+���Zx����I�(;���HT���8ۨ�lU,\J�����]���WF�����TQ���յP�:bff�,�����Zg4�e�VX���ዱ����kB�J\O>N��Y��~2�~��8��]*F��("���;��O����WBP-_":����o6��.��jom�A���~�'��yۺ��
|6"���J�����刐���]ww����������&/+���-�
�;b#���p�]�T,j�Ռa
l�l�s��`2�adD���Bi����%{���m쭿�9m�Fꠧ\Շ$5��#���
���Q�5M�y��r>�p*�����i�:kk  ��\K�L����	��[�x���Z�br���P0���,�\z�8ԝ�i�58B0:6]�i��C�V_�(G#��{�l��á~n�."�2n�T:w�:Z�,����%��
�|���ȍ���A�7�z�|q�DY��j|,��ژ�vF<]$��kFS��F�2�w� ��zlخ$�n�����<Gko�;2 �Lz�Mt�ELB�+�e���sxݐ���4[{����N�;٭Q�m�N��L�ͫ�r�=���]��[��+���W6�S
>sc��* «�(c�����Yg���#��ír�6�14'��~�פ��Lܽ�Ʋ�.�S����&��	�s3JR�S̓�U�@=��D;Q6����wW��ś����t(
�ݏ�@��Í�qo��{R&kҶ}=e���A�R�E�B&J�a�?�aI����qr�u�d)Js����3
N�LO7� )*�>y�?�!���R���9�r;Tt.Aw�hZ���GT��i�&56��]��u����%��.J����h�p�؂YDf����:���]`y}xC�������\�G�'^
�GI�fb'�����{�㖢p̰Id<u���]R+]����H����XR�1cCQ}b�S>!�#��$��Ĕ,7n�|��C<h������*�Wӏ|����+>H?��!�R&�D5U��[�77QO��b\��V4��3��b��bno�SFU��څr���"����Zq/�����ae�����bC*��C-���� � �	C��X����`1��X<�Xq[[H�KǾ(��DǮ#���+���Sx7t
{���f�ᬊ��JE�P3�'�G�U�Ǩ+ţ��M�����8لv�^�w̠�B�^�F�z.�p�`+�V�
�&l��n��{�����7�F0Δ�o7-�R����ˑ��������³J�Z�i�����X.��u�[���07�ׯc��J�c���6mU��<'�6_�:j4֙� �5 �qg���he��Ӓ�����b{��APb��W��)���� ��Ζ�Nݙ��jE=��oB�����ӡ+a�?�Vxű�C*��W�X|�l&�@��-W������Lr�`3a��5��[��b���&��};0i`l�{�q���i~~nz]ᰑ��@�<�L\O
8f�v�+��w�+��ޜ[?���+��bӋ+��1je&��Ԩ7+����O�5GDʍ8�8�V�w�ۗl|�� MI\'t�VNy�U���Vu�L�g�=�5T����Z[�,Ǎbx��q�a�*O1���Lu�5�>�A��.kb�L��g��g�,X5��S�۠��.�(ᢓD�/��T������ꍽ�C_`(Ʀ����t�e2��\6���
kTwd�[u6(�]��JD6zj����x��/ͯ�������:��.���I���Y����Q\\��%��jjj�UuyK�mÒ�����.�@�<�h
O�}Hw3I�"͚���Q�:�i�>1�4<�9#Iazzp���T�r��q5Q�P8���I��	�k�����r9�����{��@�E��%K6�9��Q/�1�I*���7y�y�mc�V��\�JT�@lC\8�)Vg��R�R���q�7�wo�����b=ѼA��[q]XS)�~��ȿ+3r�6���^�Ow���A��: ����9�k�n��Q�_�5}��9���4?+xw��s�xV�v��Cn�?�IF����[�3�U���^�����!��*{Ik���KO���	v�Dnuo.V��5�oa��o��ύ�킓S_@�{E7�W~?e��Yi-�f���]t�Օ#FѨ���/d�VTl�
�J,�4�J]�~c^��W����f����+k�2�����i����9$�{�Bpnla��Sv �ٓ�\�bt��O���yR��{����)�~1�;�&�M��o;���K���������T�A��_�	4β������O�ׅk�l�f����T�WQ6�'G��؞�2���l���"ň����'��_s��o���P�g��#(���s
<)�A�Z�x��o���~؋q�	їX��
L�1�6'�w��M������e:`�
q�|�А�����PeuuImm����D�gu�A���$�;=E̒�m�[�~�� �o�}Q��&~ff&�)1.���3G�^2#~q�'��%����)�����A�N��K���B�����2==4����@ۆwp�K�OwP$�6V��G�d�-�r��~M"���[xX����`icS[_��CE*�x^��'��җ��M���	��ӵ�s����I�_�z`nÍ��w��:��qE;2�$#q��G�A'�6R�{��<Y�b���kh��˥V����î tԦ	oU^�盢�c9��@��{J6$�쵳sXF�b9���̙ԥXLy����I/��W,N���58���{U=�$�dI�!�rJ�6��k+s�HǙ�*��H�k{���{����@��͋�؆=���L~�j���w�`S]q�v���,.�M��$܇�\�2NEF&�1~3M���7��߫��`�+��xA�ӽ������c���^�uXˑd.Tf� ��]�^��َ-���o�?�y�:(�b���3�ŝw���]�����Yq*��	�R,q)�町��+�(F�w����nVC���F�����7Q�X�6뤷V%�{��_'����:�,�����`���T�����F����_�6����/����0��*��9����1�����L.�٦��zQ�RP�W>���`�h]~�ـ>��w���.�\����5� �#�Z�݋$���AJ�ek[]����iX�^������9�ɻԉg<f���Ԣ���$Z���q�K?nU��� �1l<``}+ܘ��k��1j�]mm�?Cr)�A�t�\�mD- Pj\ʠwѼz�wF:�V��J������xbG��f
rk��<�Мa��������4p]����0�-�Ƚ�,&λtxr�/����n��Yw�an46��M`6��/�n��;6*��fȽ���S4%ڧ`lt(����L�1.��h�W��˂*o-Ũ��Ma���}p�����
��wh�t(��X\�~
����U��U0�J7&��� ��a���7��噄f�9jU`�*���L�
/ޔ��_�S=D�����'��pwT~���^�3淈 �淌#'|�Fˏa��d)�n2�O�|3�d�j������� ��1�A����r�KƵ��'�	�o, 99:��8��n�ܖ�wJJ t��0'�<װ+O�����6��љ���"	cC3��۔?-���(iC�v�Av��}q��Ş�h�cY�a�>��`s�+5aqJ#6�4[:w%NW�cH�0� nKL���'��ˡ���N���g��,O*&3:��o,�'�U�5�����*��U������7T��S�v�Q��)��Z�tQ<�˭�wNIR�����@:�I�1?�� �����}O�,Z����*�Y�K۟;�/y�ibVRӼ	�7c�g'�
���2�d���Z9k�@����G��+�(J�9��r��=S�v��)�h�'��f�ϙÈ,m^5��Oq]��hhA��k%)���9}�����L�E�L�{�5�ۗf7�!��5:�Nl�7ekZ�(���-+�W�l�u�7�,0����C}���rs�(��`kR4�.tR��4ۃ�L9�._W�}�Q�8A��o���@*������'7O&Iݹm�����U�$m��{�PKM��X����,j$Y�<��ӝ��{o��0���5c]('�뵕�~dq�ef8�0~���%B]������'�����Q�\��#���)���򌊜�`������w��A��ힵ3e��
�׷WL�������ιr�W���%�Q~�����M� �1����]���8!��ds���4�E�`�<�4-�1e�	C4�$"#1/s�ߵQ��[���Z�R;����a{��j���u%V�AW�M�{���}l�Hئ �!ek.��c��lt�LV�%�J:��g$y$�%/җ�u�K�F<U�]�I:핕��358�H����qJ��@ ��ѬQK]�Q��X�d����Bf�ǵ9�O��(c���
z�v�s�~_�ѱ^n������R��LO��:����p�q���[y����|�������Tr�d�k�ɓ��6N�-Z�I�mGg? �5��p]~Fޖf�Fݻ���.��^�Y��M���K���u���%q�z���M��5���ͺb�: �Ŋ�dwww��NO�F9�n���� ��b���82>'Ɵ�S����D���Nԝ��7R�m�L�P�e�W��n��6	�fy]�[k���V#[�~Jr�q��b�Lu�+���ߓ�B[˛ڊ�[B�t�mv����k0�K��~�"����G,��ϯ��a.��o�yOP6�\ `uO�]��{_��?�C��vN�Yr�����lBc4�IK+���|K���"�!l�P�U�矱���):^������$ ��em�!�K�w���@gAx������S�X$A t������0v"�(d��`�D�2Wg�R��庴��~�E��f�PƛF�15���bU���`Qi��j�`��xCx�H����\P��4�p*�s�������5!9���L��ҁ�{�u���S]�s�n���7
��5Mx����yS	ۯ��6&�ˍO�vVA��*|�Ś9;��f~yArZ�p#����p��Rݞ�/�D�e4r�Ц����!>����S�gR1���o���p�����Fs̔����ZTSBď�`�\�7
����Ưv&���Vұ�5b%��~x���A�������> _���vA�ou����t ����YB���60WT����󛃃[���h�0����^\p��@ .6�-Ag֞���Y��_�L8�B�����D�\$?&4O��w?|��Vľj�t`/?��*�O�:�}د��V�t�췗�=�n��[1ǡ��UX'I�D��W<��?! $&7�Ye��F3�f+E�3�\�\�{��>1���b
���0�>p~�~s��6A������I(!!���8|dn���.!��o��������a�B yW�7�G���l`s������K-y�(��/��~�'p�k'���	3�;�!��M�~k�f�F���$�wt��`��lWX)m����u�>���ۥ%A�H�@BRR�(�4K��A�'�ll�6Pim�-~ѷ�D`�9�W�3�
�p�-0Z@�Iso�����X�"��J&{c���J����R�����.�����ڀ�:~='<E�;��q$�m�s
IXx�%bۅp�����%��?�L�E�?,"�߅5��/�Vȴ Σ�'�8�;��ן�:�@�Բe:���������� �%	�<M��i$���ҝܞ:��j��}�ēh�9[>�*�y�3�B��N���xR�)�βW�{�`5���*:/^�e���,���Li���+f+^��<���.�[h}�3���ؘ$�C�;�w�A�yS�]��R;��O��]�����#��_�eYt�_`!�ן ��s;�3�`Vg=xj�	�?��h�s�@�<�NC�P�9��c'Df�vCJg�l�	2(ٮ�.>�`�}>'-V9�p�����Px�Y���hpː�R#g�î����s�퇹����m���<��,����ն�b���]Q���b�į�×���U[uߍ��@[Yѹ]m�	#m[�ѹ1�;���N�UA P�-콵�N�\�8s�����.	%�z7��o�_IF|S��s��},��0�Kq�X��{���z�z�e	���&��9_p�$u�*-zb�\%c>�*��kb��	Tϖ��oU�9��a���y%h�����֊�}𺌒tjگ��V}���ѽ)��Y.<#�w���}7��� ���g�?��Sn{�zq�&�sP�"`�� �@�pB�`?�v�����ë���>��T�����.yy��!�?�/�ng;�ik���
��$գ��}z�������K<�F]q��`
_����h�0�)�wM>���_�{=L_KS����["W���I`�P��	0�E,��#���i�M�u�����C�T]�uSbŸ�V��ʷ!9����	9Vf�S��c��?���[�p����H.�ח9<����,�/k��m�����$�2S��Jd�9q��/?��"������uB���K������Ϣ��������D��Y�|�o�t:��;<�k���~��-��c���6�,�/4���đ֤��h�8��1
4������J��1�"�\����X�����j�|+��~b �Լ0Ob���Ȉ������-��*���X�/�٨�D30_�C���ꢦ}�@�l��,�͎���ˏ�r�r�U�ƬU�0m�����U~�}�w����k�]��r�����U���K܆��؉���j�7�@�ݱ����cr���������6�qP9:b�e'�M�:���ƀ�J�`�ծ��¥7���f���%�H��-��SmfO]�S�*[����r[k� �4:�z�����[��F�~���킟9ݮ������~�}~��Uσi��H�=�,��b����ku ��=�Ɓ����C��}���88Tc���8@k�	�8��;a�/��9����SFN�`t�z���"���^������>�55�����(��~^roe+ , �����eq�m8��9�7�/���(G���G������qc�\�n�،k7��M�]�1���a���1�c��h�����u�x:��ɘ���q)i�U���8���0�v��ZW�+ ���~�9$����mۙm��AW�����f��ɣ��0���^������ԃ���Ĕ�l�ۢ�~��?wJ*�-�\�h\�������~����ޔ"@���ڷ��:��%5*��hy�h��\t�����)�W��>ܾ��Y����?>7U�������(*�L�KQ�s���Sr/d܌���I������3��|ח+��͵9	5)�xM������7�{ 2�>�����e�?�[5��:��SUU�e���fh��.''�����Z��@��y�l�ˏ���4>�7C�c��w�f�y
e�TnJu�Y�5o�����9��Ё�n��b���K/>�d�E�=��e�ȵR��������D�x���xL�@�5I�%0�>EԳ_k>�_g�ce��҄����xM��h߁7(1)i�p���ܸ�@qQׁ_�_�������V0��3wvv�ڝ��d���v��b4Ld��%�_�������!�ԟ�·$)^��g�`M>rB�/CZ��,��O��<,~�d�
�}�]H=�Y���,� �{儱��Ww
d����aU��o�y5`�����ۯg�н�'C��_'��������m��iD�o+3�P$���l��%qb����`M�@m^Q�_AوI��Ejw�J��:�YTR
jt~�u���U�˾.�'��_W��͂��9��ғ�@l�V��O7��t+��O�l��hS���iD8��} Zm؎8�, �Kj=�M�yRT��ˌ�_Q��U���3Ϝ�\\�g�} �(ܲ|�)����M�+-$T��Ic>!��n�eIj��f�K��[eh$TAE�D��K�gX�秺�i#;F�kEd�1�������*��B�~��
�?'^`I�ק%����p=f�dWו� ]��sw��Z���_�GI��(z����p#�~0�5�{l|1���q�+$�F��Gy�\�{4���]�p��3/o��wr�����
F$2���2ǩ:�"G�ʿ�+���Z�֡�M��rѩ�?�V���"Z�0�=ID�]��G�����w��;+$��g�rё��F/����G*�c��)��.���sW�<ߺWTVT��Ԍ�F?qp�#���ZT�7�I		�4ODM-�� FO���U�0�f�X���&�%((����`W�"y�H��က�����ꪇ����_oo�Kn�[>��ͽ#�wT��2v�s,���������=>k�_��H�۲�������X1E<0�?��>st+�V��a8S�d���a�E8P�TS��D�}��c���]1
Q{�|.��vLcB�#��8j�в���@ԝ\��X/D!����pu�**b��4U��b����(sn�/~r�}�޶$s����Q�m���zx�h���j[ * 	nu��C~�XϬ@#q����(�T؂Oe��p��07�`Ph{�2o0��Ӟ����kЏ�����s�[��������]� ��Tty�K:111�FI�姧]����G�ʚ��]��b�>Y�WE-�W;�,.,̪�ēP�eKR�Ht���̂b�ISe�A�q��g� 7����f��Xh��i{ܚ���o{��r&c�0���')|M������:<>��<v�9^�� ��?��nB\4B�:i�T.��8���P6����M����^<�P�v����;���B.D���K�	�7%�\4l�26�aP�Ⱍ�5^+��������#c�T�'�wb��j�">����~')�*�FR�@x������Z8W6��)qQ�fY9��X�̆R���<�뻩�o#�2��Rc(0�c��*ZZ�����cc��^����L+W�k���U��5�dL�œ�b��������{C�S���bA��?�:��'H�F�r,��G�Ы����`E`�Ja ���D�*��(v� [^�.ԍ�UT���k��D�o��3��<�6Δ��������p���$��9��D���^��ו��Hղ�t�������#n���f���Pʩ�q�ǧ�
��ozyK�jXC;M�xp9�M�`������>�����a�;k3�%kkq�n�qJ�~�1��kX�:�~珄��!h�&�>:r�a&�:�|
�&hS�\J&x�&p��^QBL�A�L]���4��|��)�#Kf�	I27����W�+�/�K��B�r��t���1��I�(�V � e���lٳ�b]�֗�em�#�������={?�*�nݷ��x��U H_�vʈ�ʘ�Tz�6^u�\�A �	)��`|�Ǥ��P�ϭ�zw��8�啺��LWX⬭�V�0IRE�UW����p�M�����b�",1��%���Q/n�:$���Ş��{��Я ��*��2�{�� @�<��y�ʐ+J��2!�y.�Ս*4��]�w�}�*���%,������#�#�(A�͋����畔䖕a�L���:�l�J	�-~��y/)IDF�����⛽��o�^U@�>�^˴y*�>5B��f�V�J9L�Q0*�CP�% )QJ&��=�mś��)%q�a����bn�㊿��X�����	�D��2��3�vM K@.	�"��ْ���F�6>�z$!��j����(�w-/�G|6U�B,�ڬ����Ǳr,̲il���x���d��L�K�T����0���g���Q���7��rm7�w�S^�qO��nb�y����qq�eqh���ĺ�iwG|�߮&�W9@�ֽfk�1�:���_M�9�����gN�����qe?b�|��}�97�9r���&6����m-��Y��kCQ�{�Abx������'�0+�����[ �����0�w̮<gx��5^b�?��{����n� Z ��X����_F�%*�\�y�>��vL\��ֽٌ��.i#�X@��n�����˖iV�E�q��FQm�!a�����%�ABR�W[�UK�:���qs��7��Ԝ`���˿Cl�R�s��	$+�ڹ�)�s���OJ�c�֔&��{cԞ%�,3�'.�Q��
���mC�e+�����	�@4��J-��� �Cw�����y����h�۾β}�/��<�Ů:qk�r�c%�ƾ�-��VQq���j�)L�Ͱ����[燽�w����?9��B�K7Ġb*�U?��� [�ח~���̫�e)Œ�Z�����߄��Lt�m�7D�W~<�f'�3�;���޾QE�'�FO� l7�?w9��uB��M��S$i4^������l{������lm�<���V���n+;�!�C0�C��ݝ�$�M��?5L��L�Y7���.k�̀�^\ �w<��F����)�/��BOZ[�_n���0�Ɗ���$i��
��&��G���b�w��f�"$J���G��p��z03�+�{{'A��_���cf��aU�r8{߷�����/_�bz�6>"*jV̘+�VjFUNBT�n���u=�V�wc ��ݓ�p�S7�:���Ǆ��wj���n��D�#�T��ƪ~a Q�d�}��sI�`�p�OGcM���(��,6�y�:�]R��>���ԝ�TއBW➵ ���!��O���e|ũoF7���I�G�	U�ࣛ;����������8;5Rߗ�L*E���F"K
�.l Рy"������e��%A�����'ҽ��*�+7��?~��?�����$�����h��|Wi}���$�ࡰM�z>��֘�y�N6�9<���0��d�G[g�3��J[�:k�x�����STf����S�%KY�O���Ma�(�60�2��	φ��~���@4>8����t �3�K!)5�ϝ^fYF|�_��a>7�QR���9�f�5��%[�F�����C�V,{r/:�WQR}㘄�Dy{r���C�#
/�QT� C���)�!�Ƕf(�;�����3�O�!�uuuǜ	�/B��,�5_�1�bh�W�:ӴS�_�����R��+���*z&�j�Ŷc����j�Ece\�T^l��˦fk ��r�n�
ͫI��E��㙊���c:��g4)�JmH\����j����C��CCX���x�<
����W'ph���y[�\����x�Ɔ��)�R���y���8��Ra/<�F)�qA�8�h��`q`}@-f}K�T�L��ƿc������`y�_��n��o0��-a"8�<�;�����u{%a&EңJ/��%��t��*ǵ~n���ρ���l���v�j���U<Λ��V���[�S�Ƴ���d(,n�b�]��t.���\�?���Kj����m;����� ��drB/dL��V� �O��2ܚ�`��ұ���SK��*�RAd��~�[��j�J.rNw�f6gfe�m*�<L�]��l�92���V$��fAґ���v�y���J�\)Y3���^�J���N���Y��\__��\��A���I�q�<)0@�C��7S��Y�;�%V�HrS 6=#�SL_8@Z�2&�p�hC�{V]�.�X:�� �..?X�� ##�WPЮ��$�L9Q�po� �
�P(Lt5*��pw�+4��qަ>|zhEE<�Z�d5h��9��H�����k�s�P�������*[�ᱽ�D�Ţ����ղ#C��WǶk�~���6{/3�����K������$����)1�v�ɋ�W���l�ϑe x0��i���_�[G�ṽw����2k�;|"s(�]�֞(S3��X�Ք4��x����%����k����n�̹/4.KI�x�߄�Mq�U?$4V���D�E�%\߀*mAA����{�la�J
)[��\k��Kn꽼��<1��ppp�j��?�2�t��!Р�������/�K<~ѣ�j�����`�C�E�
���Z��n�pxq����)>�n0�~�0}��i���_�B�!O�/�61�?]4]4���ǭ<��I��i��wp�s�ZI�|�!�Xz�6��&�>�	�[�^0��w��y����x��1�>9���R�F�� �F�����1�\��%�=Wh�>1�c��`��8�B��,8��l���ɜ3&���=Mb��M����Y���u���7�m�j[�\[z�߻���~�/��/���^��L-�-�+���Ő%#ҳW�� �4�b�OVO����AL	צ�����M@�������f>��A��v��w"�c̛����[.���YWW7o{&HV��Oj>��Ze+7j�PP��鍚@{�VۮD�#.Sp��˰ ���7K:Ȕ(���W���X�.�0C���{q�։�R}N�}�{�G��)��q�!P�Ka����*u\yϬS��a��T�B�cP���9*��>�J�ޞ�xesx�f��c8	�ɽ,!װ�3c����u�H+àO\A��;i�� ����/��|�"�л�UVǟ�U��7�A���`en����e�̈́�Z<3�~<X �]����+��7q�ccc��4�c2�ӿ�s����������b��ڃO���,��b��L��[:���x
Sb��dop0ާ����;���� PW��$�˭��lz�$Z�K���\�q��z҆����K�����j���aDit��u�1� ���4���U���Nh*)�h#�llBMbsgz��Q^�� �v�ec%���υ��DWdg����<���j��s���Q���ufe%���w�I���,��5��$>�ˎ"���hR>_��X�4ϑ3E�Ø�t��5,Q��@���Յ8�Q�a��e+kkG����<�U�$!4���yh^���ɺ>7i���3��x��R��ЄJ�*L�Y����o����{�1��-"�xE�z����C��&��׏�b�ťٺ�*���&{�	!5ܡ=��r���	R��aA����PC�^��Ќ�C�OU��,b�!|"�w�|~�)(p:C&�`B�����EY(��~�~�q~矾$�Si���%�JVTT��U��3�-cDDB��ڊgX4�qCSL�!K�Gz��1�6�#��9��^<zuAr-m��Q֍�r_�./yi���{1�B���K?K�� ť�*X_>[�ل�l�HH[:M�O���1��PI������JWKo������P�J��my��Mq�������v�.�$&K��gKD�A����л�����sh�r��;��`)d��L����߱��\�<ai�:���͂S�ݝgP���U:9��VNwLUɿ�Z\�~4�����'!���M������ڜIq��e������e�!�
�\}J��i��äi�L�	:}���@
�	'�����m�Ғv{��3Y��ݐ�"����3���+h>w����& [����ڌ�>CfQz��a�cj�2X�SՆ �%���Nώ�i_[�Ŗ�rI8�����ʽ���
�=�E��U�@zd��x�����8�3���V��{�D'�j��F9���F����A��U�᲋MUa?�9b[cw%c�Lu�e��2�o�ݯ���wt''}>�4�i�<�=�_���8����3}O�'T�-m�"�^<�2�l�Y"5 4!��ԓcfO{�[.��s���!����$]]Y�T��HWwg���i�&b �DI=��~��9g�4� 4����ޤ+�����M҉���ˏ����$<�F�Da�mrD�{�������DagC������	�$�GFFz���I1����,o�ךg���.N�:4��ۥ<��M/��=i�ׯ]�wleXp"B zU^��!�6�SZ��Vb���Q-r�اcE~1��C�˗���L/��1�r�.��aU����\�B7��*�J���|�u��@2�Q0��&��?<Ҵ(�f��s{��A3w0e��J��G��:��Lv3���{ۡ��6;���� !9^��4�����9}����J�ɠC	��.3p�Q�MR�2x�5������|
��q��3�EW}���"4W��3�c_��;4Hw�HwJwJ#�����%J���4ݥtw#��p���㮻�uϚ�8�|�yλ߽���7��kg��EAr������=���,He˕PW��=��?���#����=�VPg�VOo�E����	y6��rS(;vm�kuA�5�;��;�s7b�
�&Y��
̗ivپ�F�!�̸Y�w.X��i:�)B���%��D��Ƥ�fB�h�\��GTg�ڼ_�����Y"�^S�������2��L����~+Պ��ey�dٍ+��.����+b`C*#E��z�Ig�e�l>~@��WYl���a��GM��ٗ�0�3SKL�x�9��?���*%����tgg��>E�1�lмhy�2�v0|�j~'�O�K_�����_�kcJ�4�%?�m��Ng[ �v������Z/��D����O�A^���%��Q����c��Z:Ŭ�ˆ�*�6$��i;�����ҫ����AO"Qx��HAg+w�2~�3�\�ݩ���r�+_��4.tv�~<w�g}���Q(�m������h�ޠ���Eӱ_$�]�P�B�"�r��?`W�]{f�Gb*+�(rg �6 ]z�� P��NH���h��)�]�ѽm�r��f�ݶ鰪���k��_�ۊ�����^[!ԝ�6#�u�oNzJ�0c���F�\�$8e{>r���$�?5�i,1�5�����$��Y����~���oa<rn^p���@γ1�����L�[��R�d���(P��)���^�Q����L8{�A�頁ν�+�@&À�uy�;�D��=FӼ8pB��[,��+[�cT/��kM"��c*Ьz7N���"f�3����a�>���/(�۸%1ճHU����0[��#Gә�S%��>ٽ�$�5�%��I��E�N��3f6��f���j:�d�>��r>��}�Ӭ_^���A
G�xB�r���J�ɢ+!c�@����\���˖:g$��6�3Gp�с9?��j8��Z�����vӚ��*��t�oqeu��,�,��z�p��9W�ӱ}�b�u@Kk�p�\	mlln�#qWkmҊ�haaaO�xab��A�J�����r9q=�<���3`I��N��D'C��H�i�ٖ� ()E�p,S�XI�����u�(\�'�{Ԭ�����}�����̳GJ��h�������`'�Q���h;�ǹ��wen���$17RV��=�U%�}�^��l���!y�Z�vꣴ�	eFF��˔�@cHM|R���ް��#]tKBҌҮ�ުBw��H�M�����5"/� �9W�,��`*�Z<��܊��6�����qC�L�Wa�n�~�M�0�?��NJʙܟ'۞觲 �?�l��_6<�G��_^0�O%fhr+ʄ8wѤ��(s+:�ɗ-7`� �Z&$�f-���v�ɺ�Y2�s�T�Z�����a������a���k:̻���MG�A|��i�A&ǋPV�|�6������?t�\u����U-�G�6�f���;��}���k��T����z�b�G҉]R7�'�њ��a��'�7}G<����^Q����ބcex��TT�)��#�x$����`m?uY���!��s6�MGFg|+>�v^ϕ6���l���bP�ӧ���ϔG��=����ұp��ڰ��PW����q��zjAE���x�^���#쿜$ ���������:�j	���2���{�� ���{��.�v�rC��i��4Q�p�I�3{��P��"����V��<�h힥���hB��b^[�_� ~Ζ������F��]1}���)�]]Wb��Y�hI�؊�jvh��t]���y˶�x,i
�
�@��T+q�∾W�/�b͎l�Ȅ����j�H~�x�}c��Fn4�����U�m0���V���4��3.T����zM��F��g�6���|8rK�I�
�%ZI:����p�ti�9�|��=��A����>�f��0�*�Ȑ�J�+.�z���i�}&���������[k�k�Ş;�T� 1��GB��늿��A��lh�g������ά(J�f0 ��d���V;�w�FkhBBL�������j}z��e��o�+]4xS��5�!l�f����"�T	��-�0�SeV6�ytPVC�Q����C�mg��<o��H#ks�>3i�������PT\q�PHԝ���-/4��d�ہ�����r�!(�g�k���םP�$u�g�"����
T�����[�.�r=2����Gb����^���{�&Q<t��ix��}O�6�f��G�i�~\Ѳ]N��F�5 �~M�~�Fdp�񍢺�x�S*�߹��s�W��k��uc�a��uz|��[�F!���/��o�����F7��@%$��Ŷk�IǆXH�)�\͜�N��O7Sp/��{\>�o�4/z	&��K��T�֒�J�n@d��.A������{�K�+Q��%��'L��Z���|���S��#l���9��L�݋��fv;>�����������lBħ��$��+�p�����Ðg�'�G&�����>��	���MM�*}�K,��*�X�Њ��B��0|q�n1Dk��`Z��&��Lބ�@�q_��m�y4�Q�����V�JE��A_���kvv��'>a�NU9�Ղ+���I�{���Q�$#�.1�����S�bc�4�Q=y���f�ȶ�����៹;:����N�HŒJ�r����o�%�\p��r��P�����Jm���fq]�ݶ��p���Kivn�òܡ��e�ST#]�Od��iǀ8G��r�V��T���Q\���祤��OL�)�S(����2ф�&@�=H�4�D_�2H�8&��#��f79�u�x��<u�;6�����*�\ �dD�T�w�@#M��oyy���8{{{�%%���#lPb������}}����m���|���6������3���^	|/��F�gr�,�C-p�������&�/��2����͏�����a1����YZZ�
E*<S��uf�qͱ����0ф�����@S_��䟰T�M���T��K�"��P���e�iފ����ݶ�ŐN	+}�N��̯w�i��A*}C��Qf��v� I��Ě7kq��/1�ї��\����������y�k�S��"8��'L�G�zD��|J�i���a��-}�츝�⥧�swC��?w��>��x������"�qe��4#(ө���<� tx-|ok��`�����:P۫ޓ��<	x͞d��7|E~���t}L�y���/��KP=l�H`��<����W����^��ͅ��L��;�p\m���I�'!S�.��XO���=00�+�+YC����2U�\�����c-߰����a�U�T�TaT3!}���h
i�#�yG9�tٕT�i2I��:�
lcn�F�Y^�j�.��/J�9H@{�^ڳ�v���x��nk�zE�^�Y�Ϊ-DM- ৏��R3��YI�0z�hj��4S��'�X���T�p=��Hb��#Bl�Y�QQB����dr'@����p���7��i2�� Y^ow��+ʐe�uۋ��L҆��>��?��()� z���O����y�g�3 ��r��]���۾���V�N��W��	�X~�&J��~9�Ǝ�Y�01�k���a�#!�ct�;#��H/R���]5�{@޶}���Q�P�6둧&��6��W6��v,h�z#�Oꛜ-t���h�2K��򄘑;wI@���B<yy͌,�	���K�S���u�t������k���r6byĖy,�������-T~��p�Sq<���Ή���h�7���긲� ��9'�E�/�oV&& �=3ۘ�!�}#���-��(�{����CD�3`'�vRc�6>�rsL�K/�����$�N��4�E��+��=1*��|���?�q��,/���q���!D4٪�ui[F� ��J�Z�
lbJ\f�й��ĥ?��(f���dc����+��`
��0�
�H;m��	�1:����;V�g_��q �]`��bG�h�K<_
A�>���O�Z�:�sW@�n�S��y��Ÿ'��.3��� {X��̻w�����K~�~Y
��vU�cD=}�2��7� �C?��mkʸ[Kd��}]�����Ê�W~���$���b$���dĴ��\"!_"��O���x%=�Ïz4L$�Ne�ϓX�u������;��J{c,��V�TFrĽ+��_��,f+��m���,Y���O���!R���i^5�m��8D�a�����Zf;bJ��Gli\�V�r��(���&r�����)3���?[e�3ز	`���U�o��X�)�È)���PK��8���ѩ]�h��}\y�L�˿;�2ۓ����*����5���HOܺ���SbҀ�\�}2�@\�*vPٛ�\�QMM|·�ߜS��̸���*5�SS-��'`����h�=���*���1�>��|Y�j9��%�.h���2�:~��}dc3D8�\�� ���;�RnBh��..�8ēc��`�?>΋�R����ǹLrr2Vm��ɫ-�.��h"`�ax�Ao�����+��[ggl��?�L�lR��ͳ���a���d����f�]�Ğ�.3No�|�r4XDK�v;5����Bor�>⎶]�<˵?���z���X�>_t�L�z�����r|[7��4ܷ/��`��f�����W(���F���T	$���kFFZaQ����4�sh��ya$X�}�U��g�����Dm�փ��b���<@�V]�Lա(�n)�&����IJI����� ޾�6�j������@�"'*�Jy����櫰���q-��=0�>m8�����%   	��Ԥn��\D�y�����ThHu�+��֌�{Q� Q/�Y�%Cw��qg'8J�Ѥ	I1�8��ۄ�_6�ǣ�+�3�b�j�7�VU��;qoڭ�OǞO�*DSZ�oۡJ0G��3���[�P���λ�o�6��c���0[����JK�8dYt��AN���%�̣���LcOOX��С��%�H풚�lڛ���5��SxF@�<���U�� �;q�y|����[TTֺ+I9=;s��	

���B��+�Q�:�f���9
3�7�x�e�6mBg�����8LhW�/��n��`&YJ�aA�SVgSq�Zj���,B��hku���Ŝ���EUcI!���9~��G�؞�z�`�Q���F�$��k�U?$�~v͎�DL�;͔��Ue\�g�#v3���I�ݝ�[��� ߵ}��k�Y$N����65-����~���3���R[S[ˠ!�#���E���x�y�S�I��m�ScCl�!���"���dc�a��jB�=�\�	".�����89��eqQY��h\�'H\-;�1�R��b���?��kARs�4]�z�|.��l~0;�]�5(����J���E�!�v��*�y��I
�`�)��kZ���U	�ZoLOO��������!�EM*lcLq"���ں\��ַ�<As˭��ZQQ1��i|E�e��Q�����lu��#�ﮙ���lx�ʛ`�/�''ť����m,R%ee���Ӆ�2��F�R��;~��Q�
F���˪X/�z����Hrؘ����QүB����C�.J}9��54�wy|Y�{�����|�8?�U$��{�#v�x'�K���e��q�Y�%���փ7���̬s#L���Դ���ؤ�x ��i���	$V�o.=a�5��V��"� מ�� owuu��5;:D �r�N$�<ʁ��p�{�Z�һzB�h���%jf&�&+�H<�c��)ϋz�s;�gp?=�AG'���s���ZP��0�c�G N�f/��#e}���7R����������~HRۺ;�����6��)��}���>�����|��~����c8�`E���D������ A�K�q��O�S6��c/�9\�z8й�)VjT#K!jaAk�jr(&&�|1.�����e�@�����dδ�Ob��A�����`���f��dђ֡�s��ԛt��4�j/\���`ddd�����3`!����=�������:-��8�]Xg��.n�r����g��z���b�$���N��o7��ģ��ZZY^(f�3��?׺�QH���{(F���m��答�l���g���V���n;]"Y4,�^`��1�o&�,������m�R�wq�T(@���[�/g�Y���nE�d������v����z��~yqQN]]]OOC	+xxX�Y��/�Xlƥlŉ�^�g��-7O�$Za�>~�e�Y��.F����[R$)�ۉ=�BP��t�N��I���*c���ys����S-/4�t0KNp,f��̟��q�e#z��bcUVF�F����G�!��שTB\?ajs�u�g��-���xyݧư& ��fA�Bܹfo�4���x�lo�>1&D�1����b��X�|�0����Y����?����\$W��~�?��ۣTG/�=o�q�}7JGWx٦q&����n���o ��_��DG��T|z�a|t##�H�UODט�I����&���} s@���3?���M�jC�7�Z[Z�9<���i���s�p���+�MH�|�?�+0�� �1�i{`�;�Z��m�;*t� �}Zg���dv���=jB�&���<���3�-{i��
�UYa2S="(�������?fRv� �������hjj�z9�������-S ���a����b�t�K9�2��=M�/��'4n�Q9������{������l��ע��~y�mvh�ݠN�D�D[�H轼]gL��B��΢�&��MB_�
؆0����w��8����o�ޥ�yS��k�։E��߿�z��tBR�HSV�����3�7���3`���Ҹ6���!uj���[�P[~���yq�P������j�3n]_�����=�G ��x�m=���V/>�/��>{�U���Hd�"���7a����l�;�І�������bz{z�ϝŔ;�ߓ�IIr���S���<����P�V��K�ൗ��E����k��n��M�҇��������J���W���Ic�WӦw����ͮ�q栺&��G�)��@����'��a"�����מ���µ�s�e�w#ս�V��Yv�t��Ll�>��Kd�~*��@>V��Բ��D��)в�8̨����@<^/q�]{_���<N�;��*��Ʋ?܎4K��.&D��H���H�P��i�)���z��	�8�Ք�����ݐ�����\S���dc�VGC�Ș���<��h}�J޸�=��h%��w'
 �m\���(���z�����ב�C�{kh��;��e�����|E�6vp�+N� ������@�)VxII�?�i�؀>]��>����8�����ߨ��b�]W8d��1`|)���s�|X2�0���י}F�1�B���Xuq��7�����y#rF��*{���E�uX��"�v&������.ĩ�˃3��^�- �B����#FpwU�:vd)12�8�5�����.�\�ϡh��C��L���r]��I�,n��n��R�i����=+5�(�u�c>��'ocل�iBhe���:R�pFzSS��m���{,��;f�cӼ|��**�םҬ,HAф\�J��R�5��s{�_3xy0"��-�T����㏈�[��&X/��%�s�V�|c�����gj'a���5%�c��RV]�2�(H3��?��O�;�I<%q^�H�=`��ۯ+|��|A�|���i��uC��H �HY�U.J,��sSUzБ�L����pY`COr�WT~�=��w��B�M�`?���sX�����_�lM� �k�Pb3��p��)����}�uT�Ϝ^��w�9����D�3p a��4�6��sX��x8�9�� m�u��0��ٶ�xU��Jf����d~�e���������m�,
ԇ~7��ުkyIz�`v/����Iu��Ѭ���^Xb���c^a��i�s>�		�u�Lhm�� �����t��I2�(�:����4H��j�}��X��"uw�*X��%�Ԏ��t�(2G�|3;>9u\*gё(�Ŗ���"�I3��i��}b��_�ul����v��w�
rex[�#�[�������!���wF=	x���q�u�c��])�׎'d�q�����=��=lp�/�%����oM[�F������S8VC�d
N��}k���S[[��fC���/=Yߩ��������݉����)	qs�� Ycl���s�����z����?"ϥ��0��T[n(�[}��w�G��������|���9������Vv!]��[��f�����]���?avY�F������Q��y�l��x)<�{,� g`�jLJHHH?�54�"���xhp�����|'f����������Z��D{�l�� <6�t�z$?]��������/Ҕ��q�d����hT��������xh�G�(�gG4��aޘ�	í���~X�O`B�A#	W3�t���m�R�/�%?C<&i�h:��Zb�Ut���ﯟ�LL���u�����W/=�-'''�`U�5+:8f�^�{8f��
)��
�0|�K���ʺ'��X[ �2���)YO��ՙ"� T>.���%�L��l0��RŎ(3V�C�s�EdF�?2�Q�x��W'�.w4w�f��N�.���G��������"M�pG��/�j�$'b=��n��R�?�`��D���wO~��l�7"�4�޴�&P��.4��GA����~�Id��f�$u����x$T'�b����d��ᔩ��[L��|�g���FgW�m�R̪��XB~��=�ֿ��Y��L&R��΃f�}�V�.��'Fa����.*2!%�\�en�8�0#�KI�;��ft`�9��'��e�0��^GG2��M2�P�*ۧQ��;h(��� v�k$s����R�
e��3�wr,������ڵ��X�K�2ׂX�ouFMI�^}Z^8K_ژ�7����qg[�ֲm�8�e�,UUi���x��.?�h��wwx2(��t���5w����T�n$#D�-"�lV"<��H���|����ˡ��2�[!ݺ���0��������Yux�i�ͰL�}%�v�z�	�k�w����P����1*z2>Z���9Oh_�j�1K�v���Ȑ��njZ����(��NH�
�[����������fM��{�s�=�τo}�2FB�33b�}o7�%ڈ%?T�@́D
��M���+��E�:f�k~d_UT�=e�8�歙ך��u[����+���i|E�m�=�5뷙�Nf�Ý�q�4��c n3~+G���بNH/K�m��5���Pr&��d&�����^���KE���6���?Ɨe��D=��"!� ���̸�*��S��Pf'/�>�w��a3�O�2ԳKY�a�N�g��vB/[�>��QΖ�'1��B����2����~DE5����	y��g���Ӊ:�\���"��eiI�a�Q�
�� ���r��W�\��-���C��Ә9V�ц�l�b�Z�_/4:p����y��b�p��w�>��O�x7�������i��׹���^����+R#H���~~B�wS�F���'sV��κ����Ճz3-���8u�a=F�BC� �N�����wř��/�q؜��a_�s�nk\�Ud	C�j˶o���^���Q-Lr-�Ou�}"x
���0`���ܿ.��r�q��Ԩ�Yy���4�ə��ֆ�_Uֳ�w�VéT:���J�{goR�ʬSp�3�k�{7�+�8��ѕ/���h0��ż�zehm� LV��3::���.�:N8�I��ͮ6��@�E5^�ז%0ˎ:��M�� o��<ڃV�'��s�0jP;i��������Á���\�,�Pr�vY��6gۊ�����ۏ�u�[eA9{,�_(]]q������[չ�z���[��;�q}��/�s'_C[,����Z�䰰���P�-�;����>�>��p�����C��
�F>P(�DFF6����EL�m�N�)7�Ȳ�����1�� +=B��L�����'��ϥ�f�*���t]�a��㹑�+_\�Ä���3z�YVpK�ZC���g&++�/�|�O'�Z�_��*,*�  /ߚ��^[z �5�&&kC��4dHF84Qm�Ϛ�t
+����aG\]����AiX�h���''�A�VL�!ԷQt��%�+�)�y[�>���ӹI�n�p ?�si�+� ��.i�;-8�$ha��٭��vU�I4P"� �[i]��;q{W�:99�����\�g�w2�ힽ�`P����0�9X����_(���gٸ7i���O�Ee�һ�no�u+l�7�Ma{�t�����:oٖXN�η�8�DkP���ӡ<�w\-z"hr����v�V�W�Z?�F-�{���Кƭ���\5�N�-�{��@�ăVW�V�]Ua9a����-M70[FFF&���k��1�I��ӑ�8/���3>&�ѕ�GwML�1�aN/�:����=�"�S���^ T����`��W�% �#`�G;+O�j�_5�׭>�Ş����M��(�8�75�����E�_$�,���*�tKVP^���{?ۑ�2�aŢz�V�Lzݿ�����F�9p2=`?S��\<<]�	p|����f欥����<����+ϕ������Y��|�d��4Gt_�����[�r���]�/�&��_���3�3���\m�kԙ�~^|T���hB^82ڄ/��������~g�5�����Ӎ�O,���7>XKkER6�r��9�HHX#��ّ���t *��W��+
)�8J/8�^�}S��*����f�������c�˽�\ԭ'�ژi���-��'�Bb��wfT�ݿ!��ޙ����0(�%��׏}����+MLG&���|1dו'��ָ�������
���A�9��Ѡ{:]�눩���?#m��-���v������bi_����u�.՗�&:�At{�W�κ��|�k4�����5���{lT��iM��˦3;;4��{,��c�`BS����8_uh8&��:!Ckoo����(m��+(���X�x_e~aW�z��ROL��E�,d!Z�b��,S`�A����(a\6Tl�Wີ�GKU�&�ya~���|��k�+��m\%������KOe�,�yw��.CO���,,l}YC�?rv����Y"d#+?�o�ԋ~Mnc$�2=s�+��I���jOG@��o����V����t��O�;���fr>����lg>�sS��lpڶ��u�6����%N�����f���]�Y4�� ��}ӚF$A��\����w�+%'L�-��p�:.��7U��q�{�tzh�Gx~~�V��S��� �Қ[���-� ]>ٞ�M��N�O�o��?���.�pu0���,�_b�=E*h�}I��4�&)�(�D�����ZP�g,�z���gj�����d����劀I�~����Q~BI[QU�P�����7��i���J�mXc<0?L��E
��j���I��JO�5��AA��R;����<>a|@Z̖4�P>�W��j|�.~l����=5��ZW�OtF�\ysɉ���܋S��V<$5Ͻv����s8��a>j�tf����Ϳ�����q_G��Z'�N�'����� h��nY����r�I*4z@;C����[�>�#X?�"K�]�
�l�%���������=l����#��J9e,nݹ$�|Ԅ`V�O��e�U��h�����]�*���mP�a�1:�X�E-x���ڨcM�c��ك�ī%�5���F�,C����֖��L_qW�[����{,�lo)�x	U8g�t�{���7-�_z:��\���uuvBv��h
�fbv��z��Uz#bQ|@$��0W��Z��ǍP���fw�@�Gh]�I�g��N����ٯ��D��p�=ݜUU��~�;*�o���%1���䇫+������S��oЍ��w�JȎs��fo4�3����$1_Hn_�ݝg@��7QȻ��h��%pZ��T��s6�,i�'P~g>�l9�lQagg'l��K��qE}x5c��
,'��ٖ&D���(jd�8���
b��2̔f$��-���y������tnH ��)�U���²��6V�0��%�e�����Y�9��m��"/+C �ʁ	����?�� �Pk�v�n�!���~BQ��n�A��e�n��q��q�1�o���}X����W��`�V����\�t��'Q�t!?v���%+��w�c�W��z~�(͏�,�v�ݿ&�٬�!���t��Lz	��)(غG�R�m�MMa[ZZ�w�X����R��3�{��TFQ�t&��w���씍웝#�f(K)��燑����*߈�A�eMh�u����T_��҂6��&//i#�493Uꩋ]���wؘ����֗`��fZ�?������f6KJ�8�d��9��>�/&����7�z���,��Pʫ��c!_��"B��qϷ '�}���l%�<��Y\sw�.cL%0i��J��c�^��j*��R#`�����m�;�{�ܸL4�3��Z�K'�����f����Qw�9\Q����wRE�#�ϩ�r2B�G�u˻�ޞH@�@J�3""��*�B�x�W�T_(����Li�������+�m�/.�:����;L�]��7�������'������Hsz7D����u��:/.8�*g�O#r��|Ohk�T>M�/ۧ��600�V�`�\G��w�)�+}ep�p�'��|N��{1�^��tU�?Z��C��>�o�c�;
�?�����(�PA�m�(fB��QH>}���7J8p�ȉ�a���Peq�ޱAI];����S3qlj*�h�	96��A��x1�F^�҂WV�¦����ë
c��G�yf�P�1!g'L���p��}���*�>�*��u��>�7�����^��;[۴ڼ��o_2�>̻sa��׍M��/_$�!X���l3(��}��#�y���0�Ғt0��h�94��XD��h_(�r"��E�������ϔm�^� ���<�ӭ��48C+�_��!����wyjHA��VH�������S��Ǿ�o���R�
;+L�"�@�(�
1��{	va
v{mKj�~Iˤ~I^�w4����^ A��;ᑳ�l��A<�������r�5|w��`���'2x����I�氾�sסR6��F��4g�V�u��۠��@ �Qr�Hq����H�q�7��d<d��hiW9�K��gΩ[!*vs�>�4L]�� '/&�B�ټ������GR]]���+����73'�#|�?�������c�Ir0o��Qmv�G����Wn$3K^�3��xmbk��$��l.FTs��D�{LL�XOt#���$�(j��QЌ�,"@��Zu����^M��~�L���x��y�2�2�*�{�	o�b}?ISff�����hz`J��ik#5N�*q�����f`t��k�L:� ��-,D ��A5�>X49=��!�GB�˞�a4i�w�_�}��[-u'��0���� B�Eg���y1C+��/h^\@���b�|�8i�r�>�ö^��u������	L��cb��+>���e&�Bh���1���8}�2SV��vr,��l�F5�J�6i=�/�/� kx��w�䈟)�㠿L��Y.E����$��C�2���~VA��¦niy 8R��e� u:�/�d	�0p�̗)�#���}��xER�7Z���_i6��œ��D���o|�l�����,�%~y�������JK̗���f��b �&^�Bğ�8Ĝib ��ב�(�0�ѣ��S��a�cU�0c�wy�3���h������ʧ8ۦ&`�p�w���~
h8ԅ��`14hxQ�M�?�(��晙3&�8#�0@̎�������.�o�G��9��_�7�w�������>�.�7o5������U�۾}|��`��kXnK�akGw�W /_�����Θ�w���(���0,��N%��Z�!�隉A���LGy�!��o������m����X�a��j�����_�>���m}X?��-T�����M�����{uA0F8��ʜ��%��=�v����1o�����"�cǿ��3�:�3�\�U;"$%r=��o�n��,�����Z�W9*C<ɢ���>�����M��$���"� ���(�OrD hpB��C&�����R=�v���}x����BG��^�����e���D�.�$�pz��������p���a���C�ͯe�Yݕ�(������94�	��e!)X�t�Tj΂k�T!�P�%r�D`V�S�3��t-0�� fGq6O�J�h����
/���� ���А�Oϡٱ�;���ʹ��Q��FXE�;�G���;̄��8$(Ż���oz��m�/�;C���x��`�ԝ�Ri�k�ܹ�;��Q�� ?�䝹�}���u�&���2��'���I0�
<�:��Aa�.��;��8�yVH��g�����H�����N���X�=\�!\�^�A�mR4���e���b{�4	t��SwST��y{�r����s� ddd�[Zk�p�c� 蘜��t��J�]�B��viK�S���8�Y�)�?�k~����J�v�W��>������tT8�Ï�U�y�6�J�>�E|d{%1��<�Z��p��sj~vn.�T���_jj��(�c�a@F���	hE��	QKK;��F��S�+��2��J)���j�p�o)���!�F6]��~!�|�ڪ�h���-J�Ϡ�7'�*�n�u<z�C'އ)�j�@��
@�����6�� ŒŐ
�5�Д�A�����u��϶��?�(mb�/]9��Q㈨��Z|7� _�n:޿�����=��~o�N�+��i�?�.m�5��[L��HdV21E�J�D#q�����#X��I6|Q쀅���F���_�SU�XR�Bhj[��)�kŖ�z�h:�k�$�k�M�����{�/bX Q�BB�b��Bl[��)�_iC��2��2(�%f�U�9���(�ނ�0O�G4�?�{?9����V���Q=���Sˤ�$�0��d�����KCnˇ��R�=7��i�e��k�L�b�U��KW����V����n�-w��	�L�Dӻ�����9�У
E�.�~����.UUut$XVV��=����;O��oM����0�f��ҳB�fF�Z�l|fؚڝa�Ox���޾ͤ*���{����Fvf�����s�Ao;�N�+K� 2�� t�_ U�yj�9�����dm��-~gsB`_5rN;��;{Ѹ�xz�>wS��{�K��z�ɠ�8d�B�����O%�ӵ�{ɾ�������ި{�Voh�O��IkmEij�}-;ו����!ʹ�P�P9������" `YS�=̂�@wf͞��y�@������	�2�!涶�NN�_~Q��K�_`}�n�F�A��|�o^�	#�V�c�s��+�ˬWbz����k��*8,�|v)�v����#�wQ
����U��l���Єg�t-TV�
jP��DѠ������zuJ�:X�7�l�]`1��B|�Oo��x��U<TU�&'�c��&8��AU�_^���C�����஻8�/��CgM������6�X�'���,��L��B�{������7]B�RB�:*�]����ξ����ݶ.� V�'��p� �Wﾋ��vbE{R�V����6-]�xi�i�y��1�Dۣh�ҟ �Ɩ)��=������p��y�夘��'?~)2�ٓ	eqF--�ѩ�`��� hH�;|(���D�)N+��Xm|.��Xzv������ ��zqu����N����t�3*QG�B��B t��܃>ֽ9��G��}; ��̈́��d$?��N�-�;oF�/��v��������ptn¢�c�Z�'4�	��OM��pp���{�������k�:B��+t%u���F^�o��h���5>��Dj�Y�A�7��%(����?;P���C�� sX���7���c�O��Аm����d^�Ť~��8�ё�+-/2���z�{��(�#�g� -�7���͆�9�5���(��'3t�������
	��|�2��-?�jϭi��t_�lU�`�xm;�5i����,�f17��&�1��;�Cs��d��*��b��:^��D�J��?�Y_��q|(����oGD=�yE"���:-��U���>>]V趽�i��O���.�ށ���)3�tY��|�>���S���f-*�g�24L�����7cgo?h<+7���;X Z��pq�W�	���_Qxzy�<�6���cpcp��8�l)�Nдr���[~[.���j��ҡH|*3E�K�F}�A�$p3+л5�p���5/Zu@��|47Wq�΁�U�Zg��LMK[;��z�1�ҦOo��IjC.�&��$Gaط7���r�A�'�W�I��$�4��~rD��n���ew�v�ȶ=$�7�./��s�~�~C,n�� sy��Bو����ڍ��Ga��A���17�t������9"�9^z�5�����5hhh��i;�*ٗ1� Σf,��x*�3�����i5t�|>�b��N��lC՝q�?��eT�=_���%�Cp��$h���I���!\�Ip��w��<�����2kͬ���>u�j�]���ͪ�vo8ʷo�ĥ�E`Ai9�s��M��\0�sT���A����d<I7A��/WNJb;_��I����b����X�ش�}�
9�̶�\d-����/���PH�Z]��8'�r�Ůg�f�{30�8����0�Ae�^R4f�	��4���1���&�?��#��"���I��'���n�3Ԃ����I�>ӻ������꿱}7%��~�,Aw��5�:���u����pV�ˎ�CK�2��|O�8�i���������]Z����JRR˸."�U�I�˷N���oWG� �/��6��\[)�k��6?Eojf[���|�� �%��BB�%����Y���n�~�n�g���1="4�8r@����%]h"`�xD�VE�-a?����/�+�O���zQ���C>�H�1g��S��wy<���B�����u��Xv�2������Nr���a�#a��ݒ]}��[	���%f7
{{��6~ާ�%Q��.G
Z}ޢ����(�H��#	 f{��Za�X�\���є����QEb�������j�e�Ǫ���o\B~YA��Y��Yb��ht�(�%��L�J#
��m�K�� ���Ƙ
�*���bA�z$��E���r}������y��l qKK��K�} �'��C/v'�=��a�JjĭW�=�XD�xƲ�_5�a$:�HP'��4���Ԓ�����DOA3�m��s�`�o}��ciAe��N�&����7$�3�a�U��L�,�?�]�}�bq(��́���}���'�5Ո=�z���Kˋ'�ѕ��>?=�e���̘?{x*bF��2\I���7��G�ۏ��u����O*j�iyj}��TrE�o��ȥ�rj�I��u ���9^%"�M)<>v pX�A���R�����9_��zϏ?�w\�4d'�$��~��)؆�*ɑHD�h[K�̪YQí�<1�<�ܝ/y��`����W���t��h7e8�"gK�g`a~t�%le��$ʸz��fX�ǐL�t�`�ˀ���R(�Ă�RVV.b3�3�g�؈�c`7�����H����?x�=4Q,�9[ȹ��vx�TT�B v�uy}M��(�jy���ӆ��"�hsm��f8�|5�L��~�7n�J6����L�%�im�� ];���"2�e|�����j�������ʂC�2�<�!�6�s�/ ������@���얜-8��ws�����G�����b /_!$&��핬.7�N&E7���=L��UڽN�^X�B2q���/��7�����w�&���9�f�݁^v5�c[c�7]��k��HM�KE)��;�.w!��	|���<� X���h����<O�1����L���{<Ԉ

��	X���]�>ޟ�ɺS"���{���	�����BX	]�ڍ�2(�_\�i\�ľn�r��e���?Y�^�l���u��n�����m ݴ�,t���k����c�^jf�cț����}WF��oTZS30�6����2W����/�ŀo�SM�����1�
 �g�!�	�����H�"���=�d�E{M�.6��:B��r@=v=8 Ƅ����7ho޿@@@�J�?����̔
���9Ԇ����R�5kk��;UeS64O��f�����T1�`^~�ϴߊ��# �А�a[r���
��S;�kI����XѰ�i����Z�~I�� �uI�&��;-Յ��n}���Yo�2:�ӫ�|@09둡�OƔq��-��[�\H�O��k`���Ve���3��:E�ps�"�PdJ����*պ,���>�Q����MU�9zdE�S��^>ѭ�(hd����Ȗճ�u�K:E��ܯ4�Wd�����LM���l��vL��<e���ڿ.��yi������yZ~S_k�]��;��ykی��1�fw"���S�����`�!i�K����{b��\�#5@�mt�z3ֱ�KTkx|��@��2��A�H�����[���
?�����9��"&#cm;Zg�|wy�=-p��+�4���]]]�ړ�S�iPVI��������Ȏ���f_*:܉ �S7������U�~���n8$��_A5�H}�>u(�����Gq����h9a�1%��}܂���_^J"&������0�����8��:����=b^G�n�2��H �rr�߇k�U�Y�w�5BCՖ�7}N%�n����gg��R!��7�4���|R��41�~� ������
�n���nI	���������ji!z{��.+���ZIjf����Y�}h�{���qZ�&���0�.���i=rn��U@:��_�$�ΔĒ�-vʇ'�Ī������H�kY��f'N��q�݉\�����[��C�TZ�2'BO�:�aC��
p�����c�#-�ۡ�n��\&�	r�=h����_u�J%�lB�bRJJ���i�ǻ�T8���y���0�99�io" �-#��>���z��*w寮�^����~�l�[r\�`�f�
U��f�}?v3��r��w99ߙz�;�jN6�	�f�m�2���A��"�~OM�,-Q���K�8��p����}��{��$=I�#�[�g���j^�ʳ$�������#%nP`���d��+Q���Z��xy��h)���1�9���񗓊��.�mxߞ��������iǉ?��r�.�d�P�N���y$���ǧ�uf���T���d'D�u`���'�P ��+����Ne�"���_hMm[Mmx�#6Ы�Q�[�߭x�ϖ�d����(����"UJ��%	��I~�V�� ���K
�W��]��U��}9�l%�^c����&N���~zh��������4V�l,�&��eu��Ο��時z:V��mK��@2�um�Z�%l��XGǶ�eesY�i	1q��`�1���s�?���P"��?�(G����S�TZ��*���-GP""B6nM��'Y�y�#;5�\�� ����ʌaL��9WB���^~��"�kgbߤ����cI7	ӥTE{���/�1����R��"��׭?���ꦞ	u]a�`�����(��1��}�@r�����Т���YLuj(͂:�/PV@�w]�3Cw��H�� ���ֽ�'��������Z!O������{�M�;�RzX��Y��T��_��K���0�ny�[1K�����@��D��l��rA�%)�]�~z�>J�-cL���co��#���s���`%z����F<>�!���w�@ ����Ը���9�}�M��s�� ׯc�z��R��O���x������V������Qu��4�ļ����ݝ�&�OǸ��RR� |K�UE.!���=O�)I�B��%���0ۑl���n�|�c���+l���J�^��ˑ����/�㘾������� ��������	�􎞪͆JP�z � Q����o�|��$���y�ncKN#�ѱ��m���bO����V�~f�3�nР���s��4�Ϗ��m���'v�VV����pT��7����b��n�\Q��aqpp��$�3���#�5�~�b�k5�7M�@����}�o�Ż��[Q���G��Ū�D�Ϩ�^R��;��z�%��_�x�y��mq�lC!"��iE��X'2�ۥc���v�֔/�}�E�`�Yw&]�`�T(��ղ�3�,2�<Z�!�#~��i6�)E�<��i1�y�R�H�YO��#����H�@Uq_h���t��������aP�
����{���GZ6Ð���c9���~7��·چ�@Oz&Ko�G<!���Bt�"���>a�h/R���҃j�6���tq���aR�h�Pʳ��
w6���S>ݐɱ��5��O���0�;|�{qq
Z�%����	�iP��s*A������;�D���0�%*WC�OC�qMO�z��L$o����A��0�����E�+���n���ؒs�:�#��.�����m���P��?��w����j��\f �kοi��u�����eyZl��K)9LX��I)��閿���c��\!V�[mF����0�g`c������'vƅ-�3��dk�����>��#��p�7qeo�=��=�G#�d�,���]�f������їn
��n`���x����fz����H�.r�u �g�M�E6��%�B�r7d�O,�5ᦄ �!`3��O0RA��nq�5!�g�m� �<iۮ��]R�@�:����ϧ�3Z�g��K}�*}s���~}���ts�F /]J"O�D�+?��=3��h���D�=��O/@k�@$}KC��9	��&��>�*i /g�y-6�� �M)�W\�^�:�d�)��U�(E�4n���~������u��j�I�?����"٪�K�}���Am����
Ի��6R?���^�P0_�A�o�{2��K�]B;�'K��܀���Q���NEN{���9�G�JW&�V��<q`�K����P��P-'�?��QS����R�� �Fo�wj�� q��%�0�|��
5%��g`��}C'Q�X�r�%���R�O�߮s����OY�p�VP^]�	��g�R����Q��S|j*��09(��C-+�~�W7��}u7G\{W�X�%.w}����?�~;���h]R������5���Lk��[����u5��)$����dc���#T��z�%�t��#����*���+K�����/Ħ�;5=��C����D3�L "�h���K�kr��B��7��t"lkk�0D>+��cߏ����3�'�Զ~I��X�|�ǎN!��+��r�d �l�і��ۧ��}���FwMw����&����f���a|�'�jꤤ<w1���kO�����W_�Oq���~4���w�6�ú�:�,_����p"��X�a�?�Kql�9��RMy%�Nz?�r.=��_~Is��j�+g�G@���^m�,liy{r��OO'�����<��n�h��d�_X�!c�{�s��붵�v+�`-�o֑��C���Å�U4��7�M���O���H9ήڠ�UC5m^Ǜ�J���=h�7�n�PU��/l��_e�<~��h��7z�Q 3/-/O���ҍ�]��g�C�$�&�a��!����㕒9�lَ�tҖ�67�/����E*HF|�4r4���\�utt������6#"'�!.^��͎��:�$|�ql�v�,�4���c�mF���X�����/%���|�S/᨟��� ~359Y[��TE�E����f666�rO�,�>T^�)n�"*^�*�֔}L�>�_��y�{�|c�6[��ꛓ��,��:^�9����T/�Ѡ�gf+T>���,��2I�A���1�U2Ч����	�]g��S�0'�u�[?Q ���������H5 E���σzy�aPC�����u�,1^�}�6N%V����ۦ�ᑫrg�B\m�E�v:�ot21�\5'��1��6�F^��a$�lOC�LE-�9�0�Rw��JF�_0��񙗓�1F5�����<, oNoc���H.�q��&��;�֞�Yu|v�������&����1^yamuWc5�0��j�E%%q�G7?h�B�I�%*�N��s�Cx?�ې$S�!���2�[g�e�$�M9`H�S���ͬ��-�0�\#����X@�+bRa�I2';FV2:f���3ǄW��S�0���۱˾�7EC����Or4�B�t���qc{ͻOVb��rl�&[�����,v�S	��<������i����|-G�#/Ye��yX�@egEkԷ�Y�n�E�F�������*�V#�����Y�h��.��Gx���DSgdf^�J`N�q����s9:�X�Y~����0���"HFA���t���H�_0r�6���t޴�cm,u"%S�4\꿰�M�K%״���ϥޟ�&���.� L���F�'�ޠ�-Z�g����NT��U9�t�ɤ6�r�,B9o	F�4��E�v��u��yC�*�@�#As	��ᨉ])JLq�&`P3+���(Ff�Kj!_���@�z"+�&~:R��\1A���DŒ���my
�f,
�`�`q������O�q'����$��@���/r E_T_����Ң�;,�3�wk�Yغ�����`�QiS	\�>���"���o�D�-���g���Ok͊��,�Z5�$�ͫ`���Iv�P^0~>� ~>3�9�T,6�!��R�U��B�c��.CI�CC�E�vwf�N]O4����ET��N��ae���(}�k ?�����j�ē��(���?�~����Vf�U�Ā+J)W�y�Bf�}��9�p����ǂ?�!ѥ\Z��U�ijG���M������Y-�d�>G �����c����@�6g�)-WEc�b|�D� ��`�yG�F��3�x�U!W�,i��V1ڪ�f�T4ݿc�vV%����M��K���]K-��?���(�:n���R}jTi��
�F��� ������	�,�H:��B��~�~�l���JI�Z�
��nx�:�B���frD��r�[��J���<����.O��̵�������u�S��6�H=�h�o$��2��6!��8�<�"����O�<&��嫻x��Al�_k&w"�>[�UY~����G�	U�҂+���ܶ{I���R!���D0.��B����8CL���.�.$�qaV�VX0&(L��L���y5���L�úu�vR�Ъ�nm�į����h&b�ڷ0)/�5uT\)�Z��C�D ﾤxq�^̒u�~���)�;o��3�������(���`|R�D�^n>�+�.�q� S5��v�U��ֺo ����q|�!��2ʊ���a�Ok��})�F�$@J"�2��g$���d
C��ek^=F#�=�Z͊��vQ�~�����Mq���7���2�Q�mщ���9"zb�z��G��u�o=P�<W�9���moUs�4d����W_�YYY!5�9z'`�dU-���������5�}���	.2^]y��HX�T���Q��G������Z�W����]������FB[:���y;A#-Y�Ç����^��v++�~U�;.�G�	+'��֤)��������^��.�;�e��k[���KˆK��!��
���$0���32�E��?>�����mlm�1���3���MP|T}�`��_1ƺ,�wﻥ��2Q�/�
X����j���?R'˗)�������:��:5(�LHjr��U�YC.���w�#��+k^�t��y�tBT�G�Y�?�J�|5�1>���|wE�V����L�W��t�5��B���!3`����C�Zڬ�o�@�3��W���n�`NAA��Rq���~ݔ��N4�S]�;�3� �}��ԯlao��J�w�<�Zh;��$���7��m�W777�W,��	��OO��&��U����buqv��8�d��T;����!����ܛ��i6���:��h-XN��Q�Y1_XIp���L�'�Y�/���>��K�*��*�����	����hʯ�>����7SVsfZ�eH,�9歍��tu�$�����x��X{���/m�;����tey��/�/ �=krA��:\8��B�G�w��{[�?5�@��Ԗ��fn&�K�`L���&hjC̢Zf��
�A�?�0Q*Av3++����,��>OUlx��ߨn�鐦�����*ˬ��1.^O:�
���d�q}Y����/��]���:�����z+$*&q��Ⱅ)�^SGG�M�&bTP��g�߾�?��on�̰->��YK�]��8�6�q��-��&�uM'?H�>T9?H�A�����e?q
Qϝ��\�k���>�����Y^�gU� �
�ܯa�>�|/.ं2��^���q��b�?9���Ϧ��
��Mk��q��?<Q��S�$�z���]��/%Ƃ�j�q�mt�����-��F��s�	:jqE�/#��o�)%��3(�{�X��]i�k���ڗ�aP���4�`�i_d>#;�w�����e�����Z��P���=�4�H/&���"�;�Y՟Q�0
ᨍ钞%���e�UA�es��=5Z�Gt��J=�o�(Ji���^��TGZ�%�
2��p�����zzBU�j���Ų	�NE�"ˤ�)���Yu�LD�,%�Ֆ�_Y��-��z�VU�'x�g�qu��%�k���� ��o�a��}��ݴ����ԇ���.����T���-��:�.����ê��Ml[Gi�3,��ٳ�C�u�	&�^9İ��	�KA.&vy��wϳ������"�Q��w��9�j%/�x�&\o�3�ˋ����8��K2T�����|��Ԉ�kP4�&հ΋�&�k�E�}�_�Q_�aҷ��*S"u\�_dR�,C�P�ؾ)��ы������8��������B=�4K�}8������1� ��~º�V�_h�d.�!�k`�qhEl���΍1�<.�;�!G�6�F~���wk�8F��|�'T��o>�q]�HS Uf�B)�(iG�-��\�}�K���x�EQD���`b�&�xIe&�;��L��yЯ�%%�[�w��o�0X���}gCh���k��I�>^<�0J��h����b	{"��#�=G����;kq�-2T)���Ԧ��� 16N��fd�b�8��]����U#�����O�i���Z"$���X!�\�:��L��fZ�*l�	�ꅰ'#�P�#[����DHH�n���˔z�Kr#�m��wn`�d|���e�9��4�c��|Ѡϩ�r6��X���x���֗ �x����VH���\��W�����E����M�L+id'�\1q�I@�Ȉ|���m)���yJδ-�Yń��Z��hO��R;ц�Z����<��͂��2������'6�	�v		AȽ�І���
�X�f��FGK�EJ :A��$��Z��`,�F��K���p���x���F�-��g}���E?Gx���E93�J���.9|~  �CvZ ��.k�E�k����畖�&敊a�fGr�H��؜��i�RP]�S��ﯮu�:��`�ҵ�kn���:�)+�	@�:�bcc���ɭ�(`��@| ��
�;��Y
�#���f-��d���7J���o��-)|QC_�Tk���]�Ǚ"��?ϗ�����wlJx�?�����A�L�N%ʍ���o�VYy���qЏbxӁ���9�J+��h�=��<�ۼ��[�=!S�㨼�:b�咣��e�������/�fz��.1Y�"9�������T�mG���F{���U㰲�l[=9�ЯG�kkj�4,����b#�_)-�*$~RH��4�d��Ѹ�#)�B�����.�^,>��/�i�o�{������f�Ч�)+T�l��Q;|od�������.�
������#e�¶�m�����3��M��r��?>)i�Ɔ�U�~鬍<-v�ݴ?b��a���Cumm�ڢ��${_��!7��`"aJ�R�U�l��
ߝ��˂�
���<� ���׌L�=*Lv�7���&��L̛��O�_��x���)i �$Q2-Q1+I�(t��	��1)��N[++�]��.�UjZ�i�S��L)I���B����6����|5���9����JT888ȃd�$$p��)88�|���G�]�K���V�uD�)NJ/1����A%�c�^�y���F�{	��O�Rze�ej﯅uXO�w��V+$�@Z�kQ����6���`Z����fOv��k~B
���4~O�J	�����|��Ψ�X)]]BB
̙����fBv#iu���
5��C�=#��i�o�I��� 妚�ɩ�_��Γ�GKS���S����%ʚf������#w����D���9���i���@��8S�'F��� �ߋ]ӡ!�
��m��"a��@��7�QO��9b�~IE�0��0!���[Z�yvj�<���s>Hpcd��Al*���A�23��=c�a�v;Q�=hm��@��k��5t�×�� ~�r�Sy�]{�5��0�9"����tY�������O�И.�U'�����8�#�w
�Їv\�H�b���U����E%&��	�\8*&ym馿X������Q����R��SrI����jA�m�!�i��dih����%�t��n���������l�]�,��K-G1�ÂL1��@}y#�N�v�)W����O(&z3A�(";Z��谭���֜���p48�w����u���~�<ˢ3*���g0Y^I��L�������уS���4�(��w��<W����G"���@��f6��x`����<��8x��S��Vt�%����К��V�{�#%SR�`p �YeC� +���8��L_m��E���l��D]g}	R�#���i*�N ��Q4V�]�����n q���T;쓈�N֠ϭiσz��X������1H�Çا���n��}�w�f�5��>��=-��=aH8IYY,Vb���C��C\��������=�TM�_�Z�F�������`>|`A�,�+��9����өg��A��/���5����dYܨ߇�����IIPƭ�v�Ϳ�d��F�Ԭ*%]�(رH��:���e��)y�M��>C��'�m$�V$D'ۢ[̰'�?�U:�(̶W���N�� !�(�'.,�B^��4��z��`A�͍�N"�������#�[�صP���̶%�6-&<��o�@Δx8�.�6=^i72�1yҊ#
�=Z���ĭL����LL$�q�co8�	�����d1_��� �"/�!-?#��|�y������++�Zk`�����Λ��&��t��������k���&�6��������'A~:'�֞Ղ�����s�s�Fә�S0(D_(@��૳;�a�d9\޺0�ʚ������A=���G��J��^��"�ȗ�h�|�vǤff��|�ߡ��TY�4�io�P޴&9K�thbؚV F>f1:��YDGԎ�7�-��ﻨ���O����G�W5��~�1S��+3v�48ґFEy7<\��v���JT���:��+(� %�Ѳ����D�����5��{�K۹<�E�[ۚ��`5#O2�46��LG;1�c`�_�s�()�P�Ecn�\}k��r����;� Kٹ�[28Y�JG�v��թ�9Њ��6�����f4n�N�%���������J��Ϛ��'�}�5�;���ڒ#w�|�1I��tL
<�"�mJ��ǐ-��^����WU%��x�J̃�_�/�x�ݡ�/3]Lu�0��Z���8ss��B�T4k����])���!����7M��p��Cu,1Ūr��/�N��J+��0�������f�N�Zi#�;]�ie[�&�փ�P�jp��;�?*�>?���.�rQm.;���]g�^\P%ćR�y_�{I���{B�D�� 2Jhc-�܊��ϕ��I �X��`�>Ͽ��CW�lA8uu,�"��a���.+ .�u���"�K&�4�N6[b���;���(22���S��g�,��� *|��>>��Ԉ��IG��^�ny�J�ǳ����p,o�n��GIJ�e��_�a����n��ۻ���l�KGS���`$z��BݜY�>��Dy��9a�H$����*�uc��U�ý�3S�Ɋw�b�z��w/���:��R	ƧPxHH�-�۹��*+H��U��B�d:6IK�tw��΍�=]��tJ)��A�ڝ@.B,����R��o�����B�VW��Hy�n59FV�:�m�q�����f�n0�x�n���h���&]ĝ���5�c�g�SFS$$�KN�؄�*�,0��_K ������xf�(��a��}�K��^ qZh�U��/`g��ǻAd9���AdW��|Ua���������2�oR.�ų���U����ݵ�b�-��$|�D��Nd��&�C�$�'DPX��ݬ�|� � e��Y��JF�g@K.rO���fpr^��3�#�/�ſT�aQ.cj:ɓF�Ј�k;�Zd���`�ҧ�~��k��lz!��9g}4o���RA��Ir��f�g�~�Z�!� 5Ռ���=��Dһ�;�!Ώ�[|vA��G��_�un9!����3���V��7�`�հ�>������\�����̚���@Oݦ�n@����Q)����:ڬ��?P���)G8��Z���w1����0�̀_���[���Y����d���3��;Ϻ��v�0�' �{{VK�r+%�{��� \�9-���=W�0�� {���b@�~x�@�D�V*�����fj;��g"~�7x�D鷣�E�3�����-��?cp������TD��dg�AI���s���HZ���ޥ�]�$�ϗ �ӧ���[�«��&�5 �Vo��h#�q �}�x�j�Fo;@vm�J�����c8�����P�����/M�����X��@�� $P))w��e�M�:D 1��/(*�9���4ɪ�� nhMm�h~i��$�V�Wu��9�-�GDeR�/j�)j�{���Pi�%�����B�� Z�Mػ^�q�_='g�x=��]P���9Kܓ�W"E��.V�4�S&C��qX�!���� lg��0x^�;k��)ݨ��J�:9�C�	j�B�k�&�Up��D�^��9Y�LK��ː>��r �+*����g�,_���m,ɭ�,�%�?ߩmS&D��4�4M�W��{�����u���ч϶{䋪]���wY�j-t�:؟�o��R�|wwc�US��1�D�Z	��q��f��|e�r ��f���\��-]��B9����ն�v�rHHH!c�2{{�v����#�A�}xt���r84���1@�GW/�¾�
��&�`@��3'r����J���zs�Ӹ3z�7��;���q���*�{n!6k��,`иm�`d|�DU��2�4���Ͱ��`��w)�]W��|ɒ��� a�t��%}B2��Nm&F��r�г_q��c�#+�ct����&���P�����X��e�7*�2A������`�,�A���������Z=���SD��J����>v;Ю�s+%0a�|#�
%��H���(��o�É
���v�D�V(]��Hp�hE�*d�l��K�{�) r�#������}�vuH�� �1��:2��6DY�&���;9��]�� u;��٦�=�����I~��t=�����*�xJ������!+�Y�۽xd5:d1�R�؊�����ps�d�Z|�|*�sߎ7�.xo�$��
��ךqȝ때
	� 'Nk�Y��5�h%�$5H�D#��#���5׋�#� ���xԟ���k�v&�Y.u��Ő�e������/KLD�Ȉ����PC�8ëp�z'Iw�J�E��A�������rh�[<r����X�����֘�{�C'K��'�L����	���R=�TW7{B�"T�,>t�TT+{��i��$���L�0a����osvÉ�������U���u7�Z�EWǿ�������}&�>3���w���3"Ω�]	��h3��%k���	s��!Ӷ]��ſy?㣫�-$��M�4�}O�;jpt�O�a�,��5<bwq�5�x�P\�!�V���gQ���Q��/J?^Ku�
´�:�P�K
��**��4�l�띙�*q��Ұ��%��4�y�Dg�����7� ��N����*�� ]vC��_� ��NW���2˹��y��/�M�޺�w�l/A�:�M�BF)3@H	�����U��7 Ռ���SXyB�$�vl�s�mU�~����R��ޭ�)砾/
���5<�Tg%���["I;$e]+&~�N�Ȗ^X�SB����M���~�i_D���d��^��Z�J���!�'�D�% �sN�Sy�w#��\��9nu!�kD��#���#��x��Dxa������_)�t2��5�B�ŷ��3�P�VQ̬�1ܣ�N@ͯ=�kj\�}W�  �J B'���Qv�|�Y����`����5]e�U����m��&���b��)��	<M�8�3���̏˧�\�y��[� f��oQ�Դ����g/��Sq�
t��<�l��_���s�<��]�p�a���JӶMg�'��#���*�O:���FɊ4���5}Y����a�ͻ��?v����h�� p�0��j����"G��=��q3iҾ�I۰バd�aܦ]��kb�p蹕�b�)�ZdM�F>�hX,�ND��J����Ǳ�tn'%M}s��F\@�o\�����@�(-Vq,2ż�Eb"M�m"�>E�������8��1|ۀ��Ҝt�ӣ+ �}mi>�(B.�;�eϨ�_u�����_<O ���p�0zU�ܓ������*޷U��3�T��>���l'a����M<L�C4&�^���LB�䚎��.G��-��%���M���M`W� ��M�X��+$��8�����G�8� X=:�����9�����{�߿���b�-_P9�>п���#����	�bqc6�@t����\��V�}7G�z=����^W@=��%:6�Qn��q�Bj
�� �vlDj/�%n�f-�o3��7/����}�y�{ю�C��vs���I ��^!Hq`VEn�nrDL�Md��|�M�o�C3T��� ���,j_3Y���a>�qWr�^���!�l� �8�Ͽ�鉒�k4C�$`���h,�p-3Y�D�<϶w�A��3� ��O��o^�	���C�ѡ���@ui���OR����g X<ք山)U�Bz�i��qi�z�����Sj}���ްWJ}K!4R�~��x�#pp�Ô��v`f��i�B����|bP�#E|hf�����Sp�� �o'/�!�����{��n�"�
< |i�Xy�-%��f^�{|���i�(�vtt{��n7����gg�F?;<�ai���nO�	��OW=kSR�Xbê>�w���D�lI���B��T�V�HbS�:�n�U���GDB�lT����N��%�τ��%���NL��e�˫����~M�Oѽ}X�\�����H�	���s<f������}Q~O�ҝ�>��Ê�k���
�˵�v;;��u�T�¿-��ԬO�bS��ƪ��.s�v�hq��k�h��4�໛]��F\3(���s��w2N�5N�C'stoo�mD�~�ѝ2�%{����-F�^��f����=c��z#��PK�aW���_V=WשfOv-�5����j�ͬ����2�sUj	d��}�Y�Ure{���|���S�ڒ}�87iq�q�.<r��h��hҬ2>���u1:FP$�a�%9!���6]�W>����x5ƾ�CkC㲋Ӫ4c�����Y�IO=�!>oS���/�Es�盷ur;�=w��~8L賒����t�4�ʯxVtA��W���lC���]Bv�J�O����B�B�"�J�mm�EvA�ݮ����vu�ZZ���û��⼷�K*��҇�m�"��{|�����n�Rz��0>>���L����0���G��R|N�@>��9^�yjuw��m9�9a7�������"B�qD����ec��?B��<�$x@����S7��j�=�T�
Mk*��d�mD1�C7cl�ed}��#�A% c�^U�
�<��))�����+����R�F��e�c zC��<F�!}�O�"�fw�[/T�@ "D_7��j�z[��ތ^vc&_��-�yX	|��xx���!7BV<�XY��EJ�/�B3�O����r ��OÌ[�}Я�,+1�(�A���ݒ-ǿ��˯�j`��6�5��~�ӿ��0af��~~��1<\b?�J��Ү҇۞*D؀fg�����5my�%�r��P�M�>o9����D�ɉjF�D����-q�9/E ��ǖ-��p嚢L3�i�:��?SrT���}�n�,�����i�����z�"!�t�0��?��y۳c~���6���c�Xu��.o��k��E��25&>~ĲC[|�5�N4��ռ�����g:�]�Pl���u�͎Z��4W@����������xfd�l�z�W�8�e����|B�X�B��q��i
Ў�|�����*RЧ�2yQ��}��ě���� X��~�=���ꆐ�r�Л�*�ĿN�2��鷥�"�
��m�t��T���nl�fw���!Yvr�wt��mmu�{*��P`�ja^��d_��/���a՝8�u�nķ(�,&�0�P���3D���In	u�T'&��Yy'T�ω"�y��k����0�1J
c L��B���'%	l��|U5<M
������P�s�#�0����[��������&�HSc����(�&��{W���:8��c�4f�_C�D�����h&U$�mH�x3rNJQAc��J��@%uw�:��R�-ԩɔb���0�sJ�}F�Ǎz�h��V3�Y�Ł	�wۅ����u��nu��_�vV/��uQ�M���x�"0�N�md{=N.�[]!6�H�ٞ�|hix��Ǭ�g�&�������::�g�{ƨ�z<������np��;{<���(F�Ip��
�*����ǎ� �n�@��+���jgZ��$�R�H���c@L��x)5��{���T�/1���z;�wF����馉.�<��<?9���p�L,�c��̤�YfI�!�"��j�긨�&|�n�^J@i�xIiXB鮅��)�ERjD���$���Cb��/?��^�̙x�33�<��>��G č�:Bo:��gE��Bފj�g:|�5�dY,�ə�Qn�I��LpH��sN���0��g�4�g�v�I��Ϛ�x��<�8�ON��@ռ1��7?��])勜��iz1xd��7~��v�������b�p��ѧ�?d]��V�\̦��>��}߼�P�������Gÿ�����u�5�Ҋ�)�"�zzz{��ڽ����k�9K?������O`�AW\���!��@�-�~�	�����⥦�6~a$���l��{��j�0�M/�����G3$O�rA������ ���\�fp�ǏJ8�O�S��{�����4�V�lާ����w��]�;�g:�P\��+�3�==�M�����-�I��U�qRff�c敍DfRNΠcf\;���Z�*�!����CCèa6��2,�J�^G�}���n�w&���������6�Q�d�_���}*��
d}���W.�ͦ�}�7S�����H��EN������fbY_\Lx����$K���������⠢	�m�aV]���~����6ZZVR��Y1��˄j�x�\)--]\Z��d��
�V�Q�v���a����
�n�&��KȍiE�Ƶsv����=)�ۑ�$�Hd[n2�nwxv��R!���@\PP �Z���ZR.�� �w�������\{;��P��5��D6�^��00��r$�hR��%�Bx~4��l2	����l���͝v��k$H73���O�qs��D
)'k���6,�bX�z��)�"�9�o7ϙ�X;rU��>��6��Ȉ:�{Eëmd��pj>�"l^Ji�%�-D��?�{4<G�)�Eա��9�tףe�$5����c�, ���P��}}4�����666!4�~�p6��#t�U���6`k�I���ܖwp���d#��&v�Hc�쭺�:��3A!�NF9%���@�X�-�e<��� �0��Q��Z������׷#C��^�Sh?{$=ߨ�)&�gd,>o�����*
 ��*�^|�����jk��8S�G�ԡ��5��5Z+j����cP�\QuaaH�������X���:�A!�����|'l'
 ���ag�&M��-T���;@��0-�
�ڟ��-W�z�x��'w[��Ӝ�w������ry���Qe"0%D�̋�����4��q�ͳjMGtKa��i����%���}��3��F0�`�A�zu� �� 6������>�F��#͐Ȳ��q�F���m���locc���]t\m��@Մf��g�\ν�7Ь����C�w����u,���i�?��� ^���Ü�=H:�&]ꑷ��m�L�*!{x{�����eQ��H�pZ�IЋ�N���d�\�$^mܴar!e6(�$�Ix1�c-�(���a&�ƚ�1����C7s��"�l��F|�R��ԙ��?�]�=,��P�N�C���`q1u�DG��{}	�̝�j�JĪwh��E8ꚠ�"��J��JE�a���Y�K��O�t3�G*]�m�Y�n��kfU:FmG+��F wkrU���������#����9�K�.���f�eQ����B�+��h����dZ�`����kD��nT�_���'#��J�"��C.IIz����\��9��s�dQ"Z������*q�˳��+��\���))䃐��&?�ĬL�������;L�qF�����W۫�y�K�]�|�|����)�W��N�\�Dqz�gS�����BCЈۢT�K6�lȩ� ��rz�Jj$�~�̐��̫�7Pf��GGS���v��Rj�r�l?<����M5?�����Ɲ�#!��4�_ݓ���ܬ9\���	i�*�ȁ��S5.�Z\)+3�DLr'ąw���G���_��6b�uå@��Q�O�ܮ;�J��L��
�r���y�v³d}?��V��B���F��O�d%�N\�ߍ��M�&'����~�|GiǊ��г�R��	���@I�r8aJ
&x��j/���d]>�_k
���R;>�0ܝd^�[��~{g5�o���M<���ٝ%Af'�<�t֟ �Γ
���H[c�rwJ�CC�Gž3J�܉_�2s4��\�`S 0�N\���B�
�&��>�uu,9���WӞn�%�Ȼ�d@��n���sM
��������$?6W����{BwU\=�B�|�nc}ZR埆Yq�9�5pGVgY��y㵳�r�Ȯ��X:�Qr \�"���q2��ʖRCM�孭��۫R����&��-�V�G<�<��=�Uc��yx��54���@H�ghH2�5}��(j�^T 9�
�~��po�_P���"�gE��΍��^�m"��� e-$jЕ��d��S�.Vt�Q�-IH�����J��`}=���tT���Mq"�>	f�t}DMC��zX�-�"lh�6��J��C҉7��:��D/g���T�:	M�Y���U޼����BZZ���;X- m�����ۅ,&{ҡ���Ǒd�Чd��F��*�W���x�pP�}�}�N�}iBp��^�h|�3��G�1��66˱�
�ъ��՝���]�����fi�J���3�[������b�ܬ�2�Zg1��m�����-�#�.�z5��g��(u#��[}>�k"��.�����V`�t�av��!]T��^F�职Q�GШ��KԼX�/-�;GI���Co��akp���ՖK	�x|��ix��7���((r�����DZu�W�|[6lr�zTX��]���f-�װ�;϶�.�sZ��܆�22�5�����´����q��t��g�J��;AĂ[�}�@��n��������j�e����!m�r_��ۜ")ۃ�㊨y����X)؅hS��_b_v�N5����h��M���K�WU���o�Ȟ__YvXwG�5p�}=Άr$�`R~d����#H��+��,j�C���=�
V�R�,��=:' Ph����9Ǿ�y��j2%�O[	ZU�� @��P2�fh�5rt<i�+�F1o1���j� �#��P\rD溟��a�<��0��j�F�dK�rq����&���n��G�T�@}�D�N~~��(
�A������"{���ڝi�ǥ5OV�Ǭ�vW<�����vq�����mS++��4��Q ��nN�����b�����gii��_N�"=�1n|��M�a��n��z��<U�0�cZ���������N�o��qj��p���fP}vR_���.������W�N����Ũ�$n��mz����y�`Q�o\_�\N!�]�7�y�L@H��{�� �3��UO��/�^_��n��7���[;��f�UHr��P~����Q>���eW���K ��׏�ԟ>%�|�C�A)�8�E���&�Ī*1Zz�����A�b��ʨ�@�u�/j��AM��&��n�&�V��U��7~��lq6���v��ְ!�q�x��3����D��Y߻'l���r��>�"��p5����@�"-Чψ8ۮ��?�����3�b2{(��@ �=��IL�[�j�qM���Ȑ�j����� ���챁�{_�o{���zy�t�nt�%z��C�ɘ��n��������C�*R^k���ʔ�̱{{nk^2�xxJ��b���AAr�k���h��TCˮ�o�DI�p��"AH��f��	{W߭���ݻ���尻t��ԯ����8N>�pBo�H�����]G��Tj2�|M���(oQ�v/}�=ғ�Ŏ`�kնO�˼w/Tvȡi�N�56UĜ�3��@�3&�9��"�JJt!�W�Z���"{��=�� �HB6"9r$�_���-�Nv�&����"�{i>u��6��c% ��t_J厽��� �o��M4�5<�b|w��5%��76j{�m�C
m<�2O"��q������3��-��	v��e����t���D��I-���$�q2� e��9�1�]N��7_�vt8um�u���&&�?�y�$&V�Eɀ��,v�>�;Y	z�2O��,I�4���h�{�^퇶�-�ګ�4���̀����3�$��V�Y�	�G��o%pWc�(���NzD��U�4l�d��T�-#=�j��R�f�ݙb
�G�}�Kf�ӌ9��j��n/� �d ���5T�5�AP.�C#K����P;�ۋ;.���Q�DDp;����<�Z�OϹyUu�/ȌE�J���:Ǳ��)\��=��sJ|�r0|^R#�("K:}u�fR�����G�} s��1q
���,7���6eU�ҟB��9��tf�lU��[��������f`�kt�!��!��Q
��k�q� �y���1�*k�Є��������9��o�;]�9����xQ��ˇ�au���1�=�/.w>zKFL]d�Qܢ�%��u`y������ls��S�	ܛ{�c�
�L����x ��zȑ�υ5,[ou�B���%�~c��'����w��"��[��ܖϯ�=����Ja�G�7�~���MAޫڴ�R8��l;�+����gs̻dMC��,Rߞ�4"p H��7�ݹ_U�"_���{J�>ȹV\/���=V����h�U�~h��c�\�\|����c�9ET�甖cAGz߃s�>���4#���ɀ9��	W�_-Wx�!.��)�f���1M�ݙ��;3d�oE-��U/Ę|��l�|�`�>���9�7��h��\O�ܩ�P�I\r{�	����?d�J$x��$b��#�\S��B%��Uˍ�t^�9uv�Uu �h���d#;�-�;۵|�	Y��T��<$�_f?��@�)X4Β�2�I�����I���x^n'�t���6���eOO���-E�r���F��*�ν�,����Z��@�����I)d`��j��U`���Ӣ�T�yB�N]������	
S��v"�?9��|ugۄyґ8�#5֒��iYH��&��H ��ExF���ˏ][��[>�׬I�ˣ�J�3������C����I_�63�]
g�=¼>5��~������HQ`�Mw+���,�����t�Rj*�)2X�W��Cb�>��4���lP���ճ�r����ݳ�z���3��L�8Cِ:|��L�]F��Bg��7�i��|:ci#�Qn�9�kv�R���w����՞P�#U΁գ|����!�䦎�7���)��z����o�!�q�l�����8H��^_3�QQ��}�O����(��L	��^ц�/�h6�Qrc�T��k��sM}�����"C��sf{��0�Y�,#	�8����^fLT���?��,��uN�����f�=�K��I6�ˠ"�i�PD�[ \W
qX�>���0��U���
u�,���(̖G�h"�7���}�j�����	mQ��v�L/�'���&��Fh!EޓٝL��!���1f��#�S�G1����ŉl��W�P�ߔg!���H<��6��T86���kE�]�!�\��k��Үn>�%�H9r�wEss5��R���-��*`��H��,�Z�Z�^��4KE�j��jb�C��3/�﹔+�@kd\����u��^d�L4�.Dm- �bs�$��e-�C�o��������~)��&��7<B5|K}p%�����F5������2��X�ݘ6���k�w]�0"P4s��Vd���tv�@��=��;@�؍�q���'�)�"kAs�����p`�5��ݝ�B�,��n��+oٿ�N���yjî������+o��j��Ɵ3g%=�͔�,�\��nz����o�����j\(?)i�mp��~��|�h:wY(Ly*.�w���VI�@/���I�)p��-�/�J<��:\�"�53��rO��W��L\��e�]�T���Qt�h�jL�PM� 򳡅���b(1f��-N[ǭ�0X�D�LVtk6q��w�����No��K�tf��X�s$��r��M�|+ʷ�� `�ߐ�Gn|gFe#��#%����ZC�Ї�/��*�n_��>x��ΔR��	�~�5�6,'�`�h��u������Օ����wf�P͏㙴�B|��@�5#�r��~�pMN�@�צ��e�k�V�:�<�k����r��D&�\�UNv�5�� c�R
�DV4[��ԝ����_�6���F��#��t�"'5jb�
�%I�DA��М���߻��~(%����K��p;�G��M���#���GkG�'�l����aҼ`����N�����Џ���/���u7��󢻟�>��<=�.f�-�%p�۸1Iܜ��z��#K���&DXeW��|�+�*�ny�5ö����=��o�ј�;���Gr&�f��C�ysT�xs�nX0���\�R@�N6�`�L��#��*!M���B	�t&�~�n����;(pE ѥ
��:3����Af(�'k;���h-҂�Y\ǔ��j�����i�ǹm��p%����C&1R^�/�XP@<�˕GՓ��E!��{�Q��|\l>g� ˯�C2�rA�F�����҄��]���w�֎��.��	�P�0�i�fɅ���쓤ڼ�*_���92,��{���Z�X��y�7F�l/3ċ]g(�0P	��!�ح�]���r����Ҧ,2��ϡ�O�"YeM눺k��u��x��U��W�j�Y��'~;���U��6J��'�Ǯ�Thϕoc����佉{�%�ui�r1��>��f������������;��eS��H+*��Pl�0k"�	9[���z�X���PY��Q�������]���U����"}���q��Kc����h;��*���"�_��83JK���(̈���!�뎝}UA���lS�ڋ�=vڍ�#�2���ţ����>v��#��S 
�v��k>l�ךJʜRzu���H�+=?xb$l��m*���u>]��Mugf{��>�J���!d�_�22c'53ٞ�(�����}e�0Y�%��SW_F���^�'��}��^�l9a�P=F�Y}�!V�r,H��ؤ��ܟ'&�}��7�I�bn&�q�N�[9ItlM`���fw�IQ<��b��n��zql�Ɠ�P�1�T՞�\��[nR��o�g�i,֢�]	j�?މH��J0�%���oc�%�����x�'.���Nr�����_���g?�����+���?}�;v-dP�ո��g��\G�������/Dvk}}���,ݠ�O���e�b�I�M���G��d�������� q�����Q�%�lN�px�M<�����ag~�����=���!%��L�ގ�O���?��f�HPT|28lN���&�&���!��~|��-�������DoMȝ�
3���[��~\R���z[��
R�d�����?��FX��:�Ht<H����S.��>����w�� 6��rr�/��BÂ���(H����&)P���W<|�cs���<~�V*xHe�q%���yT\aX��ER��oJj�<QF���[��Y��U���l9%�Z3�Rf�[j��.-	���ԧG�'2���ID���B���H��mX�C7e���.!�^�=��|�e����u�$ �<R{�Z�l	�PK   �sX�Rr5�  5 /   images/ed2720bb-136d-4736-b5c1-9714f7ccc33b.png�gXSY�6@���c!��cE&�;l���ҕ�*EzO�(�t,�����
J�*5Ajh	5��Cq�yH��~|��o�./=g��ֺ�{����g�_����)�	����9}Bc��`�>q������ ��f��W]`0�S�o���a�=�3'�/yƎ�pe�00ٿ�ڴ��E�=��͏;����1SV6�[��`���9��w~�K�*�%�6׈�Ǚ#Q#�˿�Mi~?���u�Y}��!�+�~"|P���%�1[�ߊ{��}�z�|�/�?�X�~W�@z�3f����jC�?m����q�9���?h�lĻ�;x{/��YBS�"f�uF����C�<���p_�y'7|ÝWj��x���3M��#t�R��s����W&�j�0�pKb`��/{\y�T������;�g^u/��*Z�~��n��M��JH �h{�;*"�t9d
9\�fMϚ�ċ��#��.�]'o�&&E�F���MܓꝨ������8�➣�ϟ��X�g>�1��W"b�������9��p��ut"���xx�+w���ȳ��!S�|��r,�����ʫ��Fp&���B���R���!F�$�}��K���!��N�����ӷ�U�$^f*�=;�	��n�X�w��r�ܟ�@ԅ�kW��O�ީA9���D'ԋ/����W�}�H]���ǉ�3�P"n���t��j8��ܕ�l���eȔ�ћ����=��L�6b�E�h%9���Þ��3w{������1�I-�v��,?�+&Fp�g��؊z
?|��AT���{v���!�*%����زkAf��ΛsK�f��*���-��O=�BRO���'�^�Iy�y��_�1K�/�6����`nkk��1�	���Έ�8��8		��U$�1�hk��v6�M���9׆�<TI�歈4���ѹnNZRQQ�v��V�k}�T�ӥ����،����y��+��:B�JO4�4d
]\PX~m��v���ޗ�W<2w��@ʯ��E�3tJ]b��3 <BnDv�L���QVA�*?��mV��oߜ�ܤ��7iL֗��bV�������O>�A� ����ۋg�����C(�����[�I-���
�a��=[��������=FVfO������l�R�e�F����2�^l|��W��\ �N��KOx+��M|�������C�Z��n�G�������-9�C`>�:ឰ[��q�a #;�233���C�s+��0���?��M�^�VV�ec�>��
)��sޥBR��.���8�Ԥ;�����魶y�9hu����<���=)�r}�ֆL��J���M�ܹ���3�����|)����3!�1�Qi&3#cpk���C�,B��`��!Khǫ�W��\�|�}=D'D���~�i���R2�H�r��"�Qc��D ��W)Y��O	�8O��$�8Drqq:C`P>싄T��c� �H���C���J�֬��zhxh�9����Ǥ��J�$Y���t��"|�]}���A����XoI�� QG*m�^'f�;�e��/V��2��у���
^(+I�|ǿ[*�\�	�)�<l"�����x%�*���,���Xߊ^�(����}�L�'o"�M�n��[1!U�����n��*>�eQ�U�o�-C�e�K�t5:Ӵ�3R��n-�.,�+�{X�ݐ����Xh��!i��-mH�G�9�q{#���s�K_���G �+��oQR� y�P<Y�4<<��<d�2��N�ݩ1rS$�wcfg]'<J�޽��q���鷅�s���(AQ���ǰ���q�X��/�ÇoR���UmV�zh�2L�6�iF
�`[��}�f�}"�d	�@w#������}w��&s�u��?E�]�����!�Jg#XU����48�Ю��o]��~m�"C�8���o�>����f��M+�#>~~�����J��n�j6H���#�hP��F����[��|<Mo~ u��;1�Z�����r�㵮�H�C��Q�J�zb�O��4\qr
b̥6���@����[�?�U���ë���[���i��S�����C�D�W�I-��]*�ADS��q-����ܛ���ɱ�3�4
�P�F@y�o��f��i���q��*�痨i���ϟ?�	���rV{�6��b�/�A�\��&����
6�J�[�)�<tOH���t_�n���t!Js��H��;AiD�*ixk�C6!y��ґ��j;�H�A���C�i�WIt�B���h;�+�W�#�#��<�;U%�^پ}�p�������KM���������l�M�gS���/���@jR��뮃tE���rvl9��Ձ�;w�<2���J�Z������} �I8�}���a���Jp�Uapz�y�S
�YgK���]Y;�I���U!�~� $��b�������$~u"��L�(�QM���@*^ �@%�|���VO�E�{q�K�&q�peUU�.1+�eH��ׯ�S[^�A����4a0��Ѷ�3Isss��I�����n�U��L��dû�O�K`
0�[~��Ͻ������Z\����3�J�C��ի߄cy^�a���5hp�v/$�һ���o1����3>~S̽4Kv�kHK��<����u�*��K{A��#U�,q�A��F�p_��/_�<b��)��yqG���l*7��!S9�|�3��M�Syyy��١�6y�Z�l�aY-p�9��(�c�Pu/P���a����o���:>�Y)5��+�����Ӭwi����{Q��7'v��:+
�`��e��I����h;���q���bR���ה8��h�8��Zx�2#;�@{VR�|L�TJ���ϰ��;�`����/�,(ƓwNӅe���.�������zw'��F�@�]����&�п�E��K��bYk�m�=o$~�v����Z���|	̙_4(l��]P�gzf(�5O��]sp�<A��_+޿`y��mb[�Ļ@�H������1?�Y��xC�T�8I�{����j���V|jii��"p�Am-����`�73�e�M�5Gr�k��)װC�(q�AZ(���IF��X?�����ڦ���ߛ�znF��|�T�jm)/݅(��oPRk�ǹR�)��-�.�m.�N[��0
����3�}�3��SS�S���sR������������Ġ��x...�q|暰|�m���b��� i�@�ZE�$��T\�}m&�յ~`�/��؎��[K��HB�����6I)O����[a� �fW�9X֥��?�K-�0��(voKB�C�fa�R�¢"�Q����X4-��/�AFs&d������Oi,N�����q0vA�[S�A7@��������p����T�Յ�'>��<�%����	�5G����@�^��簠�Ck��R�ხ{qϩ/�&��ri��A��A����o��Z��A�����e���t��U�Ty7}]"�d���%E�S$�%�� ��ڦ2{ %pC��y��d�ɓt��x�q .��L0�sw���>�I��ܥ!��2���s_�{����Z���!y
��c��d��v�TO!�(#�?~���q�ѭI�[�6�L�ي��x�[�2���fп�)�y��(|*ۼohx8�A�{k��B�H�3 ���ݢ��^>mJ-���n*�O�����!	u �&�8�ꪑQ�nkF3�Oy��bV��|���w)��]!$^W��_�ے�x�Sm�����ʈw:h[�q��-�d���4�c�ǌ+��XI>v6 s�>	��S�!��,?��B��'� 'ȴ�@W�3����?¨W�"ˎ-a3�6^��i/��+M��O ߟ�,��^��A`�&@{�d���]/��*$�����z$D<*y��Y�]ւӭH(qy#�)8'M�`&s�,��s8����ȐY�?텽�cz�@�T�'�PO?�N���da肝��Ŵ����SS]t�L���,�_u�ЏԳ����e������rM��f�!"����L�~dd�{��ٱ�լ�N- �gK�Ր�$v?|���ݔߤJmVUn�9���T�j٘	�7�n���c��~�[x=�����P���0{�g\�niS{$<�e��|Vv0~L�����Q���]^ᯥ��:�Ra�T��5��2x�"n���9�LU�cuʦ�eQR��(��?�J]ȗ8B��Q��]mZe�nVQ�F��ֺNj7�c�!��,$�4��H��ߕ�0òw�2{&�)	Ԏ�`��T�J7D��������A���(���G��HH��f�ڙ�/*DxvԘ� 7G���B`�w�^ñ#��ުQ�QȞ1S�=Ȇ��.������t�t����|���)��2��݈� ��8�8oEi!ߞ�q~c��g����:�EJl�}���~I
w{���٬����F5�E�T���ʐ:8dԬW*�c�j���j{�3��'��M�j`�cY!e`��|��L����y��ל���Z��U���VnOCc�:��p~����4hֳV�@��{��Mf��& :��h�Ε��B║a������O#x<��O�w���TZ�������p(yf�l�P�X϶��`���A�3U�I ��:NX;���W�k���f�̓��Ntip��(�/��<���S-(�
��>`�N����R\xo��US�T_���d����FPd<�-��zA������e�Dv�O�N>�/���iS����O?�aV[
�Oŗ��DY��Y�_6�1���O�<�E��ւ��ؠ2�[���4ogI�ߖW3Q4U�O�;�-�����b�t��Hp��r��Q3RQ�3
�]9虙�%Z��*p��3�B��S�
��@����!aaR�q�0K�&_��f�׳}��|!V�K��M���1�K��!�HR�VL�f��̯�(&�ίS�eJG����JFNJ�R'=x\U��M<n$�9��ms��N��N<ם��S$�Rh-aI��xb[���:�+�� �za�����ê��*���i�ղ�x-f��w��t��MX�$�`�L�Թ*?�(wJ�,R���s;$�e�qr������
Y�^�s��Y����G�=�]"���2e�]�j��������z��.��@��p�l&��SC����q�
M���V�g��I��� �^�E��jF����#[aV�*Z^�l��8��v&}�I��	�� Z&p�f��L�\��̖��7m�h^O5Ͱ�Ɨ���M�Sq�G���Ŭ� y:4�ߘ���En7�������FIkf�l�<������\�;�Bv]��[������G7|^���J`g�.	K�ӟD��8q�x���T�-��w+:��-+K̊��D �J�J�|��0�@ufP�,�?ڈO(\�,��Zȧ�c�gT��ʖ��^��[w�a�K�{dvB��u��E�Y�O�X��\Di�:�n:w�ɗ��ʞ���֖����O��H�/���
�|y�b?��J�hp��Hh�@?����,��>ګJrQ5�7;H�w����9.'S��hs��1g�"T(�q/�Ka#�e�I�֬@��@� �ݫ���n2ȇ&A%��v��]��f~�i-ٞ?�d����x˱)����G�����D�9T�i2U��l��9�Ւ��^ \3m�4�'�7=�2��\�R^���6Z�,o�*9P���1���Hq���y�^�d3_D�'Ee�kQ��㚜�.���:��v��8�M����Vh�B��R�M)���;�U�W���u�9���]�l�=g�IɎXD/�Ӽ[Xi�"�DX����5G�\�!s��K��:@�$�fޢ�Σv`��y�!rӋl�{c��o�t�c2+1m[ޑ 'I�U-�k��6���wM����iR1�гFUI�MXC��5P��N3Q �}>/U���X4K��K��	�h��&�� ��v뢀ڲ��@�]�Y8��0)��-f�Z�V�����E#i��&g�{_�]Y��Rq�z�{l"����!�d����ʈ�~c	�i���oIO��`e�Yy2�ɪ�n7n����̳_�
?O�T��5(7��?�2��X��E�ٌ�a��]���93� oS��(���ń!)�̞��u���Cm���%V
:v���&=��%7����'y `f�1�z[j��e�}FscЛ��M}�����V\��Դ������d���˚&%f�ӑ���a䲎H��b��w.�̯�F�$�q�$�yϔuQ��b(4��C��dU"��
�b��R�����sr�q��V��7��?W'���s�ϟ�'Q��Bc�bckU��fkkCV��u��wx��XA`:���Q5����gEbM)?�"�&]¼��]]��PVmE_��i&Eh�n�"a[V���'%�/zU	yD���I�CIn�\YG����Ls	�49{Gc{h�E��2��(��n����x�����!�5���.��s{/��n���p"cϪ��͐~����C��
B���<?��~�kW�x���ny=\+�r�(zxM}s�CP:�ϛ�������KK��2��b!�O9ҏ�p-�AξQ͹��|t���j�<�tF�q ?�.q����a-�sJT������kB�͟g�}��K��A��[�3���J�
H5,����M�=J��4�$N\��L����rT�w������zj��2�)�r�/u���eg7�u�1��ng��\7�`U	'|+%[#�
aD�]W�,#���K C�;09�~k^�����>Lc��H�n���ޙj�������Q��1�EV��7	y�Hl��x�W�i$�}x��՚�$����TeÊ/��M�!K�n�:ơ���"�
���Jm��#�1�~�p�@�b��cR�X�X8��._ҡ|։Y&�% ��|k������lǄ{��};Zm���疨��YV���x%`ɘ�f��BI˞r�,��/Jξ̤TӆX���e��q"T���B��u���[��o���D���Es���~V��k�ۦ@��>���Di�����	G��bl\���j�J�[픙�
�04�I�k���~��hX���x�|�i�ϒ�V	U��Ɂ`B0Y��X���Q��h���	%3��5�w�>57E9����j��B��S�cs��0T\t�P����˪|{=D�3�LҖ��c�0vZ{�߽!>i�8QLX��s�S[0�VH�����z���?knn�E��ץ�9�;��$�o�c�I����9�5��G��xצ3yx�z��������#y�Ǿ�y�n����kQr0+\������,���=�@9�z����_��r�l�6W��2?�ӻ0	W��ߪ�3}�***��y�w`|x���Ws�������hj�æo���\�:�����A!�SLm��;,BcmF�.]��!�/p>�dԚ?�#M��S��'�T���a��(O�g%{�'�S����U^���q蹅P9TsS53����ؒ���=b+�0�n�#T�$�*U�Q����Ȯv�n��ǜ)��Kh��r���P�����ٷ,��U�4n0Q,�	"=�_����&�������Z�U�a�3���-��_�og���3! �ǻQ���x���*w�?m+��=��v��҄�R�_d���Z'�2��q��T��m0ٝ�OJ�|���\�퓇"�4!�V@�-~���8ʅ*K��v�m�:�fl�7����6�PZ��|:2
G�I�.��Jrݚ�#Z�#��H��a������i�q�N-��z��e�$X�)�r_K�W�@�"�dz੎�����?�O�>W%�n��+�WL��=��q����%���Zʻ�BY��M?��ϙ�ϯ�O��m���t`J���p4��a�*�7ә�#�ݞ�<��1>�F�ULY�<�(+�� W.G��4��񚩓i�����=L�Z��287E'�Fhow/M�صkׇ=>`z4H�
A�/k�����X��i��#��b&#�,�Ͼ��-S�������~V���}6P�U�4(�w�ﺥz��֐sZs��֗��]!�%� �rrru��+P��	To[A�����\Z=�[A�D	�b�uW���(�6�O��md֋x����lմ��a�g�� $dp!r`wS$_����P*ݔ=.��?���y�w��w=�8��O
�ɩf�w�9����|��#Z#�Iw�k����m���J�I�-D�>(9M����Ip�S^��T�irz<�A�g�� <���_eJ�ٿi+�B`2��?��{����EgQR�l(�?��I_{�#VI�Xu4?P�奙	U��,���
��x,�d�<b���K�ӡ��D���1��;|ϻ�E�|����J������N��>smF�=-P�iKjvl�ó�>���G��4�q�̏S������ts2j��{Ks��N߉μ���~��
ٚ0�7"���+��o~�΋����^^���:��=��p��pyQ����^�ޢ��,�e��0Gi�]���N��� �_��M��&LG�D�;�4�`^�P�Y������h�[8���$��tx�2���YB���ԍ��f��U��<`�xt1��$ߣ?<i?�)�Xtn.~�7^c*�;N�Ñ)��Ս#�@P5~�6�X~���h�h�3b[��i����!RH�ZPB�{����lu��T�l�^C���R��9��+s��o��hYA�`�`��
:��}5��5G���C^7��J~�ی�(�ݞ^�>Ѕ%Ш���\q_/���`
9�. ��&�Wρr+Lq��o�މCS�Ķo��j�x��*#���a˥_�M��¤���/�fef!=�C��/sI��s�G{���s�s��{#���[a]?J�.��$l�a=�o��_����afg;����P>�4�1��g�Q	�]�ʳ�����F�{�8��`gg��Oȉ�,\0���Rv���wg����K�j�!D����-α��2Q��vg'!�������g�|�Iw�]w�[����7�|v��>c���\�f������h��Oފ�Ut���gNK[%(?y}ՙ�(�9aWCs�>h4-[J{�Sm�U�}N��f\{����p����	���a��L@h��j�uT��-'�W��,�y$��*���_��.S���x�lykq���d�b�X�4�V�?�'DF���|xA���c���H{�� �:�kb�"���{�[y^��;	��zXݬ�h_H�f����?�(�+vظ?��ך���Dn|��m���b��JRrE����4���S�������A�|�Ҭ��#2����T������*+�E۫f&^��
B�XVr�m\�L�*ѿ ay6%���K�bUg{�Vqn�^��QVfT�Zs&��9z�[gU�����é��c���S�J����
jw�uJ=�-Sfjt�}��~"�M�w�0�S�r��X�r�t���U����\5]�aJ��){TY��oN�n".`�+4p7e]��!$�����0���3��$���}bm��EϪtU`vF�.Wn���9ӎV��`�;{�﯅�?P��
��^]��4x��T#�>�L�U�c]��o�w&	�G*z�A�I�B�����bWt�XO8��9�,?��*WMU�Ȓ��'߾F�z�{U�N�����A����s��۸ڹW�Y@��jy��*m���d��������YXC�d�v�Bs�r7B���:b@���}��I"��?-���Mޟz��,���ݱc[q!��󷽃��A��&K�:~�^y��0��zT��cx�&�<a�i%�+qc�.�m�-e��|<	b֕�@yDAg�
X�_~OqM��p�t�N��c?���_�����!�eW����̯_�[���lpX��n��Y� +�z7E؝U�*�V�ʷk�Lh�7��:�E�&���"x+�&b��T%U�Rbx-��Br�?�p_���K��,$�|@���1�0F�=�Χlا�y�/��Q�g��5���d*�~���O�J:�ޥ�ث��S���ga���4�#���� �J�]�*	�����gj�1e~�;���e�����P-�������NE���ϟ�"8q�Z���
q��##���F�C�y��T�8��"D���Kw�����ذ��b{��O۷9|[8s,u�[۔	�P�Vib����Z;�;?um;��B!A���=#Y�*7�0c�E�2���{��d&�&գ����Y٭l��F�<C4Ԃ�!�gt9�׻|@���K�{�|�>nZ���FZ�ު�<��M����S������HN|���S:ZZ�����J��D�m�������X��%��Zh�(-��[� �$�,L��q��a�Eno�'M�A����r%�/_�Pa�����X��,���14�z�L��_	3�
GBc�9�}�2���S���؉y䠗��/0P'��YS�y�@�΋��W�����b��qc0�*>
R�3n��S�W���%?�{�o��	�p`��|dlaa��V�Ԭ�)E��t��_]��P(-hڊr��S��7.��i^�*9�:%�2��N�"nmSn�58躻����ܺ����.&�-�Țz@�e�^Nl�=vâuv6ׄ�S���	����n�;��ϲ��I�����3����O,~�r�"�#�ڮ��N`��}�I����8�*<u�L���U7�S^�j-���9a�2�A�����si�Ж�T%�jֵW��
��������֛lWf��9�T#����%�$���za��)֊OG�\�h끌n�>�r4M���W�׻5�c�l��u[���w>�}-����=(GX¤O�������W��ڜ������<�S��ڌ|���Z�����#�B#o�e������v�k��7S��|]XȂ�%�,R2H��r�@��^[���l�� T�����n���b��U�y�7����O�q�
�׷�+q��aD�w��^��C�w-�	��9�X��§4�����s6L�&v����[Aj�u0�w�eV	��ʆ�.��X0d8/FV��,�<��L��E�.w}�ڜ,f�k�!fM1�_�܃�2��Ҋ�fQ��t�5��d�ن�s2��.T�5M
4�m� �6�RP��Ջ{��llR����ŗ>n��� ��;���f���-�1��K������|�y1�(�����z�31�S���1b}��|�@�����V`���ֺ��`�KG�o�@(�X�F�I�U�Y�)F��F<��`BX�j.Xq��>�B��f��=�<��Ԋ�_@����i�L�uK��6���p�]ߝs��՛��7�x��i�!'�RjJx��%����Zg�2&��.g������VffZ���}lBB��_oaw�4�^xg�Tb��Eh�I���E�Ů&���cZ���C�i��\��+R��+��p�����h�����i�}�J�Z��C~a�D�����R�N��A�����Χ4�=,,,:������]^���1e����D�v�ι����=�α���%�����`;�=��V��5C�V�m�oo�Wi��ko�f%CW� `�P�B�r(���I�o�a�ݿ>g�"0|�s��d��Fd[W���V.m/�]�wh4Rt��R�����A��ެ�r��l�߯�U3-a	�'�B����RSS���������}��uQ�^���cc&���ס�4 .�.Y֝w�����(X�!���L�5�����Ֆنd��w]
 ��?��f���,t���R ��}=/+�Ɖ3#��I	����k/����q�Y���Vݜ�5��X�D�RN��|g����|�_�'k���1K�F0�zi)���i�ӻ����J��xv�eO��M���[ <�S���!�M�ϸ�f��)�M�����=+oy�}�$���9#���γ,^�]ap3�1�ݔQ&�t�q�_>�: 6%L%f��<#�c U���\��`#��CkA�lV�x̲8��%7������"�/��mϦ%�հ������}�.���\� 0d3����'?tp�%P�hk�=��7[K�S���,��O�R��RpO�
����� ��˥�|~9X���;;��$�����R9H���z�{@;B�\����<���P�up�O� _�,��v�Sܻ�&��5��LL�fH�n�� \#�)���y#��n�@���gIY�z1��|I_���ye�h�}(ZǾ�w����y˯#D��H#E�A�&�%z�k��''�l�2歐2�	��&���-8ǒ�Jg��Kc�~a�c5
�o1k�7���!����%��?js�*�n�����I/[āMD#��۷?]y��~Lk�D��q7Z�R��$q�׷Ma�@pM@��U�����!���xJ�~���,��;j���:�����PM��MS8k� ����ۅV��Y��x8qm��E*FN� �(d� p�h��vG4�P���J��S�Rq���yUx���UV��Y0�r�`�~�5>h�\L� �~��� �1��5H�A���h��J�P[��\����L�B��3�+4ӱg�o�+���d\hKt`I���~q�z�u55�e��-��8�J �����:V"���?ȍA&��2�v��i/6��Mh�E�pU ��_9��do�i�Un<�n��	��؈� n��*����V�L<�B�G���NǗ�=��[��v��Պ�!;���p�:�Pٟ�P(x�l��K�7<�����i�
0���:�֞�}�{���h�7G_�l�Hg��?�dE��Ç��6o;��qs�k%�Uj��Jom}~�-�]ɱ��69%ki���º��Ɵ�.z1�(�_Uç���>�F�Z�W�#��T�G�UXqa�Ǩ�����͠�r=�8FxT"YZZ
�n������?&������Y=�A��	9��던��:�ʬ��/ �:�q߰�5;ui��g���5w�����&��UI���w|�"�n�&u?|��,���)++KV��5��v��g�{+�(��a��[�M��r����I�_���CP����M��|��"�3UC!�$v�^i�5��7.v�(�SI�c<�����$���rb�A��w7Re5`hi�`|1��O��V^�pl\��Õs)�n@R���:��<��B�QD�̪K�?mt�G�k�oq���65��C�vJ6p���+�x :;8+[mr��C�3P$<B�_	��r�MD�Jha39a/C �[�b���
敞�$�*@�v�nn��bC�}�������s����8�Ř���<Z��q�R�]݃�� E��脘A��d1æ�G������8�W�U9В��vv(���Q�@RI/d�w����>m���Mp�$��֦0�_e�1�Yx�jk)=r�ު���[�J#�Bk��ur?�Ņ�Y=IT�'�`C7�s�]||U���[u�hk�T��ֆ�g�c"���Zn"���[�0`j�/2Z+_��uE8�fx�&+@H��d'��u��M�y�����8#�z�N��SM���'�L��E���0_ ��Q�3I;���Ҟ]�ګ���,���U�χ�T�V��ŋ9V7�s�W-4���w>��	���L�Nq���-�1*�k��614x�B@*z�hY�`;�j �砉�4� �Y4��U"����NtHKéu�o��i"�?v0RCr1��)q�{�ެѱ�b��.���2%U�3�0�#��f����5M.���S� �v�}�.Ũ_��_�E���B���� �W�h,͛U#;t�xW�> '���nD���V.���jj���_�EQJ>|���ʜ�
(��|\v��2H�'�2�PV�0&�f`KO3��s�K綗����A^����_CϦ�N>�Ry��>-[m��nݚ2��Qz�	��/��E|",��:T�	���}(�|q�$}��f��U����aЁ�<��	��gϞ�F���1��,d{� P�ak����B�`/�8�"��o��������:V�� h�d<Њ~���8�zl�"�ZLh0�e�Mo����{ȈW EDGE-����������>}�F��J��E0[�ѐ��w�tGH���)[K�i=��p;
J�~6���#A<Zɱ!��~��6��Br�fC����G��<Zꘓ��@�?�͐)#F�7g����S�r��� Lʒ2�r2P�	I8n�����N5�E�O�%
���D(�=#sm��%h��O���ww>!�9�Jg�h<�9�YU��Q����-����m�>pW���,M�bt2)�����T�AVV$��I"���H��y�� �����~'�NWd~\B-����A
c�.p��onbԤJ`˯�6��ʮT��`�ʊ����nm�׽ks;r�Uc�wQȝ��eQ�R�^� �a��@mZ�Ǐ22 ���f�4%�����9���s.Dg,�IjW=�498B��|gy��/gv����}�%$iuׄĻw�@Ƽc���O��#�v�*¹w|�)���O8�|�2**���^���� ��9L2	����s�'ԗb�[������L ��t���m�Ɋ[�;~S��E�h���!�}�����JY�Pk�z�/����Y[D)g8��t�0jJ���a���B�<��#9�]�~�2���q��G��U�gQN��~���I
P����V�s��=�h�b`��Z-�*��'�)�0p暫��;1��P���gc&w�����k�������p��Y9<�g��ۆ�i$ZOo%�� ٩:))	�a��(���;�Èn6~��C_m����Nw��Y��8�����!�&��]�G$$d��F>�cM�pd{��^F�W����5�zԞ�cd�>̞Ԁ�y1�e���P���Ǐ�N�ǭ՜@�3@�R(���|5r�W\96�����>��;g@�����b���z��.Z�����!�J#hR���^:1i��ō����kA$g׫H��YD6�
��p�D��=*�ZD^��N'�0�ݲ[�`�_�Ɂ����6o%wtt@ (j{�����KX�{ 1�f�V&_�hG���ȩ�m�]�~�c�0[�Mr���������Z��r��i���_��vHLc���/|!z�1��+�1!R�S�1�M�
x�`q��<�������h���j��l���uQ@+:�ʛf|Ĺs�V��������[��ϝ@U��:�YP�M�m�������P�pR	����C��*�%?�m���AKG��0N|-�;8wlHj�[8q�mm2��� 	JII�mLUKL�l�al�>6"(ʹ��M���\�`h�Q���-��C@+1̀����.f���)KM���:P;0�e � *}I2����9`��n����xP��Y�\��:r�c���	���.��<9��M�
���0��얕��cW���՝s gmሥ���6���-���� 1���V"�/�mY���_�Í@�&�w<U��ܳ�/���b�3c{"a�7n$��Crઐ����tƞ��'+��1������O�lW�v���q�P54G�CƁz�B�>��1����a�o"�m��,��
�BJ�N�Z��JS���|�T<Dֆ�:�'$<�μ�{7tl�wz\Mۅ�Nw������5cD�J�Jb�62� `�f�ՠ���J�*�2��R��m�f��Ӷ:)�2.��s�	�D�=� �OA�?PO�6ܰE�I	�O�t�f���w<F����e�e=J{�`	��2�geiY=7�V��{��V����SV��y�ӌY�_�|95���5�4���{3��x�N�6���!�#5j{@%ܭ�³!)����5u^��wE�~�+_��������C�9��9}��J�(�z�S�����q���*�j�W���\�#X�;��˿�l}w?4�}� A�nSt>5">{#Ѻz+y,�xr�����,ݏQR�KHDf�C~������n������n�-y���F�&�����ˮ%�����daR��ųsO@�	���\���_�8_4A��0L����!ن����E�����? e�=�{b#�=X������P!���ǰ��,��I�ٿ]��XT�fgg?�T�<��a�ʠ� �.}Y�r�6��R[������CI �z�^=/=�������h��$���߭첲x?�#�ːWz�lT�,���y^v��(���\���SyI��9�ak�-�4W5���G,d@����Es��'�y�ůQ��ړ��@��p�N�&w�~.-�=a��.ʊ�&`&.u�쇈f�+���(�?~��U�Y�t�@;IF�����UǾ�e��I8�L�Hܦӈ����n.55�p���oXƀZ����2�:��܌
p�=W��o���I����𫃱܁	3sm��X���IVsgY��cS�R72g���j0� �O�p�]��ҫ�]XRR�g�iQT0Fc�����Hmmm�3dee�v���+`ԓ���쾬���|O`�"�"��^ۼ�/����LJ�v1o\�����������ԕ�'|� Uo3]�¯�@��ެY�.+˥�E �lލ}w���	�[��}�&��+����/�ۀ������I�=s��K��%f���<op˵k}$��>2��+C��v�c����i�BKY��R����>��	�9����8N�F5��8�?Ź�(6Ѭ�$x ���˱�
�>�XˣtJ?|��7�����J�^)Ֆ �ĉ���G�1������CI54��	q�������������B���o%�8�,T
:�S^@�t|f���8��w(V��Q��D\my �9�R��ح������k�OX����hK5���Β?1j�l�j]&��Kr�0�����v���ZĊQ���'4��8��=t�����2�L�ؼ�ƂN�tڤ5ϫ��o�{,f}�~�LW�Z˩G�:Tol�q�w*��+��tm�ݓ�Qۛ�������Sǜ�n;������|�ϯ�"�|������5) �gP�|�C�F�ǳ�V��Ro	�pDso�L���ZaR��!�ύ��P�/�_0�=�-�'�MY{z�|h�7�
��J[v;o�b=z�n��|`僉I�^�-������$�Z��A+�g��12t:G&�ƿx�@!϶U�v23�:�e��-Ӆn�'�l�l����jR/k�� �G�Yv�uX�w��<L��[�+�j�vT;��Pw׫܀%�Lv�B %X����ɏ6�	�`۱��r�����㡉����Wr�o@NV��~޲��|9��|I�u��Kw��rͅk!؁y�@�;�D�9qO��x�]_О���ej�>��^�f��Ce�Y��uZ�Y�N�z�~ {�1��D�!�m��OT�:�0�-�O}�:��`�*+�](���
�ﾔU{�a|�t���:�w����)g�oD������U(Z�5Q�����Ui��)?��G��k�~� !`;Q���F�K��d&�YAb�Ԗ��ă8Q���_�MD�2�X�}�՗�4`6{�ܤ�{x�A� �x�fkи��K_�fW5��'�_tI�y��i?�p�J�?ҁ=wJܺi�7ϳ�[sz2P,�U	`*a�@���	�8�<�pb�e颃������+�/�й���ZS�G�^�z�vb^�t�_��`߼���eq�ѳ+�/ج6��,�@����p����}���"a>�I5/�X��W���M�;�}��Y�1I���1�Ţ�vp>�7O<�Ϧ��1�ژi0��z���?��G���������c�l�/��G�����S��vڟ�⎯����Q��������9d���D^;�J�������|������<�o�kZ&�������_�/��K7�6B)�A[�/h讠����@�P���}��g�J- �^�B�6~͜�P�X�`9C�i���q3p��'þ�	e&�xb��2�߱37�p�Qt����كI�Џh�?e�j���Mm���ل���I_<�`�3saoV�h�e{�ɼ��]-O-W�����հ�0	ߝeb���vU	_>�]�2��8YL��:Z�G�gD�w'�� �c�o<�G�`a�u�xV���n�cYhe��s��r�:ߕ�|t3�וo:���U�wa���d~o�-���.ly���gWT��z.ݷ���6%��Lɇ|o��°)*3���Gc�iP9װ��#S	�2���V&QJ���Ut��kv`�[�����2ye����
�>q�>frYn3a�7���ٵgΖ$�sjM�)��2�u�늹����bK���yE�Y�-M*��^�*-�����k�/w����G���?_\�j��W�9�+#�k^s�:��K�Ŏ������#�]o��wP�e�����x����H��H�
]��u�k�|���#(�2N3 ��0�������Ҡ�����L��{�x���oܒ�rJ%���J5e��TR)�b�(��3�E%�i�u*E*[�)�mB�uƖ���e�>�g�,Α~�����������i�������z_�}���G���)��d���$10h���|�мM��v��9A!��Q�i���(V�7�^��ϣvYN�<��mڸ	!��s��4�.�	E�\<�dA��^H8�o�%�$P;۾Џ�OP��2L_�Oh.L���DJ{��c-���m)�+��f�)l���\�/k=��&P�P�W_aV��F~��K_�N(��´P�˸7�A����&)Y����6 �(��ͫ ��H�}��
ӹm2,�Y��9��H�}M`E ?TeZ(b��h������J�s)H�������p�b��X:p1�b�S˯\8��w��"	`�&ȸ2�q˧�o��P���Q�7�!�
�jQ�B����J?��B�N���ݤ�ϖ&�����X��/D[��y����:��ꍖ� �,�҇);%��%8`�;�����g�>}I�`�'9����N�ǀT���C�|�%��i2��@2m��3�ˎ S�f���&��G�B�	]I���k���mOd���S��3>�~��b�5���oTo�^8%S-����Ya�ԫ����D(2�~�
`������7���@I�G�Y�6}��`%��V*Ӟ�h>�(�=��P�N1�	_�A�ΐ����g�,L��]`��S��s|򣊸yH�eqA ���S;��~!�a�����29��0k�Zim�Ef���S�4 ��%����%~ZP$�b��T`��~5VZ�o�O|Ԏ��*0hC   ��ڝS̾�`q��hq�{K;���~�wp~�wp�o�'i�_�|�w����������������������������������������������������{��m
���s%�k�~Y���5�?���HCW!E���p�Q^4B6��������uGV~�@Q[<kUf�4G�3��s��6��iD�O~}�B���C�VJ7�H�bx��+P6�Sc#��C9�ъ(̋�Lg�t�h��FЇײ��^�����J�ݏa��\�Ջ�I$K�������TJg8��� ��=]9rY��^��x�@��N6���2Dxh����t�bΡ��v��xy�I�"Ngxe3��z�57�ч���>V��q���_?�41.����M��o�_���DD]V�tȶ���m$R_#c��¿l}bA �Y:���,�k��5���7��S��mo��(���5J��Y�U9�yb�*JR2�͜�,�p�~����س�dϽ�L�`��;HV�)L���SD=L�)u�\z���Ǯ�La_�H��%�ӑ�TZ��|)UPĥ�6w	��wiQ2.w���f|��X���$;��^��p�z�h'�?Xjϴ���D|�	�j�~~m��pL�a>���jė>�{��d��]3� ��|�6ᐇUX�2�9������-ԑD�S.��&c�B�43��GOM��̡w9�y��.P�p_�2)v�~��rťe���1�h����S��_<�߸�B�	��zǇ�rG�́�m�Xť��TN�E��q��D�$��R;��<2������	y���]7���K+m��# ~�5Ц�����%��>��[f�[w]W��~6k�s�O��n:S0_=�����N�2;'�˲�\���a�5��Hx|6��3��;+OmN�B�s yu>X�.1'j�]^|�ΰޯ,��8�����4�<�s�c�nw��(�ۺ�t� ���H���>-�4�L�sZ�I^������m�u�v��y�4���үc��^��x�na7g�sr8��T�w���������#5U:#vS�q�v��fAL���J�	� ���#6HN���m��ə�ϫNڕ�6��<}�mO;�_�����"���W���ե��h�p��٬�i�N0K��Oy�U(^
ao��h���k�|���T��ې-Kt���r����u���M��iYa���Æ�v�����X�Y����jrS�W��7̦��<

_���_�s��D�Y͆w ͜Μ���K�&S�!��۸L�{�i�����L�a��]���;V���	sl�=��4�u�9��Qng��2�����6�X�ι6�~
9Z?��j�ŚAt*�����6"���J��0XQ�c��'����������"���c�]gƻHb��ױo5O���o�5h�I�OIh�0*�����ϡ-<�~��	��2�o7t�$�nz��P�����EȊ��Lu����S#=�a{�j����L.1x%�J�����cǸ�z�j��>���1n���>p�&�UGU�~)�s���ʄ�u�Hq��M�@8����w��7uk1Z[ʵ��818 FY彌2��s�������j.�"u[[ͦA�%.�+�G@�;�+^���)������"O��рI��3\x=,��~5u��t�*DW�ϑ�=/��t�(�]����E׳��CJ�'�׃�c}L��ȿ"��3��ׇ����<�ZVH�ͪv_HvjŎ�*����I��Tck�}�� R��H��"7�qe`��x��S-�?�$:�a�Y������橫_�X�1ӶZ�g�OA�� ���9=�b}�Ž����ӿ��8~3`L�>�[A�0��e,���렞n���4�|C`��7.c�����4gNU.����b�V@5���%��?8�!S��$�@�D����~�Z��������^[P�$���Ϗ�o�w�G�ȫ�7�\~lԥ����/3�"|E�(�����K��@=� �׆�u�����=3�3'(��BE��)�d�m�S 6$�Ћ�M)# ����v�G�	_���:3��<_	q1k�_��8��P���#���S0���z��:J�j#�P�f�]$��r�ـ���ˡܠRfTZ'�_Dz�'v_��?�+���o�o̎��9�<*�˰/�B�uʸ���t:�H�V�i�FZR~p.hi��k�d�9�[����e�EA�ňA�p*\s���ݰ5�|�V5�J��K�|�8����"��#��B�Ǜ���a�4BsGoP�����"��_J�vm�@���N^-ř������<<T��}|�*˂^�@�9���vA>��ee�r�ELtF�fN|���Q& ��:��,�ǿ�DA~S ���Q�+��iw�ŉ���9�s}Į9%	s��]<l���� �B�E��/��$��*�q�-�9��a�� �ĥ��?T�@Wd&�����-�z!����X�chҙڄz�E�5@Ĥ�}p��ȋR����@
w�b�`웒�j�e�17�S��4��p��wegHF-f����*�@��o 5��@���`�*�o˻~x�n��5d�]�/d�.���i�X��ߣ���"
���jIWM;��K�O\ ���k*�T�K�sj:�p�,�%1v0R!�\�h��c�%��!�-�(mW�o��?A_SHṞ]���)�٥�/:>G�RP����rۆ6��=:|���x�U뵽h�jʫ��d��R4��ޗ�r��w�d4����Rr�;�zqQ�h���ה���T���Y5V��g&�=���qB�)��)|�i�j��8�Z�У���I�j �G�k/��v��ig6H��`�"3J��<��s�z݂��K���Ik�Z�I-=��,����]�!�����íq���`Y��F��Y�z}�ǽ���m�8O�gX�y�k���wf٠�=�II�,?�3
X\��˹�����H��$;tȰR^�vט�7!bbF�m=����囲�x@=o�	b#f�s�/+/ۖ����YC���E�w@�-"�*D��IǍ�і�>����6���qc7���Y���}�	�m��9���)���(D�5T��ܿ��6(�sT.�yB���ΩjY��~���#ƙ��Wp_5Yb��O��x�bL�������m�v7y)�; -�E���t��=��bEE{hi�
�]hDl�c%@��
D��1p��>����;cđ�M}��H}��'OL��~���AtGp���. ��w��{�\���)��(�b�����X���t<�������4��uF���%{�M�4�4}���>�M�:I +my��L�w_]g���f(,���ݏ�KNNb4�B��zg�a	���[�KS�/�)�
,����h��o�S�����������:w�Z�Y�ET3�n�YKl@!ˇ9��/)Z�gݺ9��\���E[�����:���"B81��AS�H�CN�vD��V��gsKqN�Rȋýge�:2��N�_����9�H�*4����Zc��$���$�69[�^h��÷a(�>�dN����O�!��"�g�a�+n�,Zn$�e_Vۦ^�v�A'�o��i��_�[z]�Tq�|�O����.U�~��z���e"��-w�}E�q*�'�J�_��2Rl�ðq�B��GU�sΒ|�$���
�a�(���iU����e���A�,�L��/<��c��ayJ"��J��/3Н�i�3T��]��8ǘ1LF��]�w��3'�H����PA�@"�ɬ���51�'֥TX:v%Kq=��ڵ-�B���$;l��&U1&�2�qx�������M���"=.���p*.]�	�bw
�$�jċڧ���<%7UqtB�;��»�@�R�츽-;KQ5T�hw1��VIy�8�-�c(F��_��2H:�Ŧ¸��dp�l�$�7"�I�W���/�d�-���^wc	(���ަ�1�n-A�^���A���o��f��!9omKC0�ӆ/�a���.F3UC���\�U���i�)ͧf�U�\�iZ����I�g�p�]��Lݼ;.����ʣ�T1�������	����4�� ��!���z�9�%�5��0/$�R*Y#-�e�����F4�BP}s��~�?5jԾ��5Y�U��M�LuOdl�&�a�*��x��O���T�:m[��j�~�J�e(=K��g�i�\P���h��z��g�d&�s�&U��hH޽E���?yaQ��P���[q�-��� (ǜ�?�������n��XzME�{u�J�ؠI9��1	�����D��>���Ɏ��NB�N-�0c��x���ƒc6�*���| ���j� w������n-P6�G���
ɣ�O��8�ml�a@i��Q����ī���^B/�)�9YG[Ǹ�;Y2��m^�ɦ�'Ҫ݃�N@ �TV�l'�'"2C��uM�Y :�m�<����3���sQӂ�r�C�<�q1�`o���0l�5��{�k�VFJ��b(�5�����[�yy��< \)�v/��'�pLǆkiDnҙ���ܳ��(j� U�ޒݓ��&��jS�q�T0�<&��nq{��΋�Ĕ��W�B���e�L/F}���,	2�Xk��v���������L�9Uw"��Δ��n�J���.g��b}�|H@X�B�Nُ&����(�u���-���;�hB��iZ�9������⥖l�/`�GU������v�����e!s��*��H�H��/Fsr����T'EF0 �*�j�;���Q^qO��ф
��ײ�"6���{�K�§���������WxA�"je ,O��Ս8q����|N3�I|1�s��l�o�2�|���v����;Ыb+];�n���;��®�;�
tl���9����{u�j{s��\�397�004�p���:#r-+6{/�ŌL]V��!�^_��Q��m~���:\�2jpR�{��Qo��L[�i; ���u�@�0�g��=�.hF�?ba����P��CuQ�.J�������g�%H�yM�@��:ř��o�/!md�p8)Q�������*3�/%��yۤh!�s�y%�/���y;sNB�㬉�<`�W���-%����� �y��F�+���z�G����@�Yo"i	�.�����
Ԕ��S$�<����/";.�rކo���ګ�{j�X�Y�1)�J���g���(��+�洭�u�'b�:L#��X������Q|��h)ë�9��Ԫ��2/,K�;Կ-H��/���%px�J����w�5��:K��'W��&��X���N��g�	������N�����):)�褫d�F ��<ɸ���`�AKE&��:ܗNNm	o��}����������.���k���r�W�R��������p�A����$�p�.��\f�Z�r��|D�w�(��'����4Ru.#5�;ʤ�Y�O�|Ǌ�:n��z+��ͅ��#��]�;G�]���Q<�qɺ3㷘��a�쥕�=łt�2����?�mݝ�	y�QZ�oa�7��7!=SB�{Y�6�]��1�N��h��ӂ���dj�s�2�,F|f��ݐq��:.�~/��z�����VP�ʹ�:#�M�_�Iu�D3�4�����3�(��:D�n��f�n��)f��!��e
�����Qǯ�-���`���8jf�50����d��t�I8�b����(����ʥ9�P�)mݮ���o9��:25�P��xT����Lk�7�nÕ��`P����'�.MOs�
y���0���P���R_H1�HD������w��^�Bby�=C�����"偒���"Zշ-�����Hsu��I�@I�/$~�PV��sؠ��m ;�B�~N�W�s/^�I�����c܊���ͥT�%E�{�ݓ�	K������.m$����+�D�%ԝ�7p�(�����e*TAG�%T�B�,Q��K��ė*��>��R=��Mä�z��p}�Uw���pk��6oi!o6���t0*|�0����72�v˻P�豑��qd
)���:w�A6�Ie8
�	��d��W�?j�&DC��=���S�D	��(6��X�����̱D�,t^IM�@�&�sq�4m]vn�$q���3��>-����%��0ﺕ(<94X
Cqؚ�*^[4�1B��?_���(�,���{��Hɮ!�`�)N [�}:�o9(�~�丨�f���j���;l\sN��Ŝ�'wʍd]�utRG��W�@e�&jw��� �o�Ȓ�p�\E(��C$���X0�%���k�.(\-�°#�d�Z��W�D��L%���|p�rH�V�׺@z�9��IC=��q��R�9ւ'�w�gC� ˢ��kϱ#4��Ӏw���R	9 ���AsK��8��~��p"��^�r~��&�G�����J*�y����c�biِ�.��6.zՀl�9���L}S��zGvG��f���㨨Y=���)�=8P;Tҳi��������f��Hk�R�#<��.��8�~;+�ь{�XdC��E�bV�I��2���=���^~�E��[`�q�.�G{��Nr�>Ms7a�6�Y�=���4Ur�f�Qn<�h>��`�!������!#�92��VI�>��u�*'�_/D��m�����A`�f
����5a���힡4cƫ�0e��;-�y��{?�B�8�҉���x2��.@�\{�������~�g������>w���\�k�9\F~�E'B�:6����T�_&d*�sZ�p�t��C
����M��!?))�;���}M��	���/�Mw����ٗwiѼ��[�1Ka�6�C����{7��ן�ߧ����>ZIH[jp|�x����p�E����ҳ,�C0wh���'�c{>}Ȼ���������m����"�sE��&��R�q@�8� �gԖ]b��+����U�x�mu��K[G	0���1�A
G��"�dA)>м^��&��Rb��(�ҭ�#l�Ad8qe�j���c����='�%�h>
�y�J�5��@�f#��̡��/m��WΏ5��ug�.�o�UC��Bԉp������Yz�Y��c�/JU�����r�u�Z�����>���x7���X��ŏ��qW��P��3��E#�4���0^g8Ҏ��Ҽct��Ls�E�)�h,��j���ewe�'>�=���?���w%�*�C�'�x%ځ{�ۛ�b̧?�b��X�DV(,����<S��zW�i�46�0�M\��o��D�>�e��33�����o�y��e2�f�W�����R���q�鐎!���M�^e:wWV,�l}{�w&������գc�{�aJ�{���VH� �)0�繯�`O��_4zNZI�?N'иi ��� Z�����!>�ɰ���:L�M������ûs�x���2�����<�1��"?�C_+�"�2\���Ow�-ǹ�0��̡���0E�V[@��ǘ��ߓ5�)�|!��У���&YT�@�X�%�-��-��d/o�*lx϶p@k�l*�e��/o �Xo���B|0w&>X�Ğ��y�b�0�#	X�����v���G�NM k�i@Й�QI֘�X�O����
��4�Qݍ�\����S�x%~"2 �C��U/�<b�Rǥ-�/�7����_%{ջjX~��3'މ��*>���/���%��mg���k'|3�k��d��(qs�H��T��縨d�e��&���T S*�����6E����j�/�� ]���������?��N-���Ŏ����-&n@�U.)4ShI�w���Q�D�+O@��
���6lQk�;y?�r�QCn�ܾ�*�����ȶE*��=�߹d�t�m������$�Ћ�G��+��x��(M��8���]�Ǯ�)E����Q�Gح��#@��_2����yY�}�RL�7x��,��q��I�yH^_z�iA�eJ�e��L���D�������>��oK^�X�Y�"\x�I�5�glEwe�ͅ��)B�]U3g�%�B:s#���|���e %,����vձ�p;�0 �T�y��@EU?������3)v��V��4�C�V�@�L�	��7�I~����奬އV��ND���fe�$
��Id��M6��[v{�2]�eH=����e�L�:a"�e��qQ)p�7
卫�>����/1��1V�Ά�Z���)�ÿ?N���k�ȶ�.$S���+�i�=|�rʜ�N��ܑ�X���f��%�O�'�y���D��e�
�c�2A�E�Ih���Rs��lM�"�����RsE�!*`Lվُ"+�����c"���aA2��==�q/����U��2n�\�{U��9?�q;�����V��������ʊ���9w�_v������ʒ�~
���{�oi�?�F�z88�E҆�	� ��q�4n�36�q�h�`�10�.?��L+����~/7M����@DD��A�����Cs�KY/����2u��@��V��'����8��J����l��"=��h,��JG��#�hȂ��/�ؖAM4�a�#�#��j�(��D9RM ��1I��$�.���1�Q?M؟^$�����o"#p~���p����u��!i$K�X�O!�RX*�=�'.�)�R��#��;84�L��`�۷x��^XaSH�Ta���DT7٭Ӧ� ItD[�~�fagط�����K+5P�e��R�-�=a<���Q�D�$��	��
kl��v?y�����y�SZ�ea�;���-�ha�v��.�x����G�#�-�4�`��y��J�n0�o�H�Ⱥ+jD���[��5��(����cc�A={A���:���HKD<N8�IͿ�,�c
�L��|!;9�����C2_i3k׵u�L�B�ք�NIe]۝�2�KYk�K!�+���7��^߆b'Y����tCfdA�!9����� C��=�	i����joGp{n���<�#��솣(Z��w�a|:`���k�~�5���%���j�Q�hn�b�mD���d����DF�f�bD���>�>����`��6�2�>��!) �Aݏ�����~J�zV37>0�4�DnyOV��<�6q0��观^l=�3��v�Md�����(�f��D��<^��pi9��Lj�w�	O_��?�}��y-�^%p�ڋT���H�G�������}�q��a7���`�NH���_��
f M��Հ&|����b�p����+}6���]Z�m�,3t�{���9��&�0��ɂ1��D.� �H���`<'�N������U�Xd����s~Ặ�2�C�� egJ/),EI��.�l.4���"9��FH	����Q�=�<�
qY��H�ߩ��<���[ۭ�kW�R�o�I�r���E�������F��k���=�q���t���0��	��7��#�#�f��x`���_
��([M��ss 0�=3����q/�;;Z��~.�� XU�|Ax�?]�G�塹��f�w2�0��ć ���A�(�&h�9�H>�x�>m�JMT1���޸vM�gH�`�J����?���BY<K�ё���ĴIÜ�m��;z���泏}L\��SI�]�Ď��FD�����o?���Ə!H^i��'�^#��=�\�����V���t��V��t���*ZH���*����*e7���e0���˴�r�?z�]��!��D��Mz��V�*��<N�^�4�9Tƥ�O.aR
��*�A�hI� �=,
#� �r������m�h�n����6Hi�����w�7��|��Ț�oonn�<�E�������z�^x��-Ýek{3��޽령Rn)K��(C�Z3��N}�u���q���_ļ���2˅�L*���b�x?�̬��#�1x�z
ű�F���b��g^}ɈZ���Q�{1��Q�ⳮ�9����N؊����Q�	GG������#���%ƿ��~���[��$��p����
�09��l���A�1m�y�o@�Y��������"����;_�-e�KL���1>��ړ� `���Z�v';F������7�����kV�A��9��PdR���`�Am��ɲNN6�Nn�����Ci�L�k�a�=t�Ui����w��=�����T�֖�-lQ %���L���A��|��Kq%r	�g�sr�NB>����K�I�DSɠ'A2��/l�w���v�6�8}�y�Fy4//O�Vw}pp��Gy�k��i	EWG�����`�F۟c_�`V�54p���`8�����8����J�'V	�E�������{��@��`䜩>�=��>�Op�\WEY��qሻ�cV�z��a��~Ŭ�2��"~[p����J]�"����x�dZ�<~��Q�o!��#��f/�,�R�҉DU�,�9*)+k�s��l�p8�>���p<�������:�杔ɗB�L%���/���!-�x-����R	."9��}}?w�NK�Q.\�����䇬���j���\�����
|�E�F����脪f��2�/��W�X����5��.=_F���c� i�=���64��٩/0ht�1�������8Y�w�ߧ����
7��z��}[F�z:�C�Ο9Ӌ\"�]~��-n��,q��fgeg���<��ݚ�X��ny��gч��蟞�=qB/vGttt�c?��0�A8q�SN^�W�}��+�KVVV~o����g��}|����zj09�Y͈L ��T��<)n���׼�u��C�>��yk������uf�`j i|a��tt?��`煍����+++�h D
_���s���G�LM�������*'2MQ�����Q���&D�=��J�9���'�Ffgee�w�V�9X���>��h����4m("藰+J^�|G�L�e�P�'�_����eP�[�U5ǚh�O���W�ÿ�,����u䘋�t���&k�ȃ�� ʖ��j��/~a8~�/V�����?HJ����M3:�|�� �����lL�Dΐ��s�?i����B�����_�ߢR�`a��2�A�v¤�b�U��V]��zig�qI�n��u]
GU���s��j�ɑ���8e��3m��u��*`�Ƕ*}f�ۛ���ɕn:d�|����9��Cr���1Z�ϟ�9��9�&d��2��7W�k�����Nt@�*��Q"���p``�/t����RcS��&��C��`�B2�d����G/.my^P�����`©����쯥�p�Z�
�R�=&zIkruPgO��֦c��H�B�����d��lȉZ+����П5�	E��rY �>��/w&B��
��� Ͻ��a1�l��S�r����	��g��W=KK^�t�DC'�����/_�{�^�Vk�J9��zȌ[�⒙P�D���v��W���x�Ģv2�k����R��;�!% �nX�Ӥ�/��_�τM��M~���mt�T]<^swy$���p�e���>�2h�.�?��j�����._:���L���^��
��bu�;lY~�������*lpM�>����\���+SI.��72{&���r��4U��+l���>�M!��.���w~m�VU�H���HHpb�e�?3�溇�,n<H�Z�����L$+��q��_����Ҳ ^a}o���H}�.�+E�_C�oY
�B���P�BavC��Wk���s���UNٯ��I����_`(�h�i z������7&:��V`w@���do�H�����慨¯�3�x�#�J�v-\��4�M��oi�Ǯ0������t�[ղ����Ė9�*Şw�{%����u����gWݩ{����Y�|BR�b����"�._I������gϞ�6\UVV�績�����[�B���������`a�Zn~�Ⱥ�a1Jf?VՍ$�]�� ����nXM��tｻ�>}b���7�H�0�k��H7i[�� o��7�2�OJ�-M���O"��o6�JO�l���S��B��TH:>KM�e��z˰�"��'0+��g�u�㷡P1`��m����k�[���B|Ѕ4��O�n�"��j� � v�����.@��7e⽓�Zi� �J���jwru΀��=���aȍ?I�\kn^�g�X���g�ee�K�w�hW=Jg菒B�Q��ل����M̉��&��{�_�����{_�*�:��TU�G��:}�g�I�n;�ߴ?W@����n�YC
&~z�a�^��:g�#�[r�/@���q^{k?E�͊�M��|��n'��^�%rU^]ũ(��t���`w�z�����n>�O�5(��@�����5�:��w�#�"5��C����L��la���-j�&3�[ FA��X+U�)�s=�*6��`�%8И��U����7�J�VΨ�}K�L��;��4s`S��@�T��y���j�@κ���yU��8qv��
�S,`��+�)�J���>�t�k�+�9����v!��SRRR���x�ۧm�s��g��6r�k���h�`��[[[S�q���N���S������}O�Be#HZ1ۜ����@ྡྷ��e{;���C��1���/�����G~��|�?�\�����8�c�̳� ���747;�S(Y$8W}\�1򐼱M���Tf�MM�н���?#3�y�4-��ׯ__P��*��s������r(���������@�Bc䪩�*����� o���9��@���5b��.��1I�Z1-Wr��'��-��Ϡ������s���QC�*�Y��UG�&�a�	N����N�y��U�Ï�{��Y<ӒY�?xz��7��S����p�Tt�����@:�k�`7+Jn`�J�a�W7W�c=�U9iͣ9́Y������{�p�C>�7���`�B!����6���X��̮��!�_���I��1���������8�8;k`���a ����m���Z*�GG��b[[�m��������|��w��SO���� �9"�FLG����s*�o�����k���GH�S�sw�x<���&3:��SY��zj���@
R�b��4ȧ�-�[��bT�Y	*����o1t���@X���=UH~�k5G��^��m��� �Z��s��\s��"q�Q
/��݁����;M��bʁ$��;�KG��|����&l)��啕������;��w���c4��nQ�r=�� �a�w����TǴ��A�"fe-��Ao�������oA���<��T|j^��W����D�x�7)��i�Z�2�>i�%?㪾�~���bm2�H'-w���V�(_wj�9���]�ozNk�~���u'\6�-1p)>�K�`b-P�j�P6$=F�=�V�/��}��ԞZ���ϟ�h�S|�~��3�:�����rR�6
8��;rqs�����{gX���G9* hm�����v��BP@Ab���ޱ���f���L!�tf�	��s#�P�x^]4�n�����+gd��g�Z_��v�K�Ә@�k�;��C�ڣ�㴳�3��tO%r6�P���xk���qq"|�1N��|����/���Z)��+ŕ_�Q�Im3bK���\Yed��L6�y�!������|�7�\)�(����nG�L�}XS!�EDFTX��R����)v;gd�_�<�������nzv6e�,�@r{d>�譓g�^] �l��(.��SI`j�����e���4���7>�8O�x�?[W��g�猩�.�h�dw���O9�ŋ�<�ܡu����x^oՌ�^��[,�e�����0#�:)imu�Hў��tB�����8�Wq�JN=:%���x��K3&��r5�6�N�R��:�s�Sp���Q��L\΅����5������wl���w3rG��6(c��W�Ő��Ҡ��*�f��6w��u�b�٠KQs�:t��.m�&�Z.+N���t"�n7��ߏ=���e���L���?���1?KI�~��O /T(���qž���ԻSR��-��7����u�=>��ΈP��G�ֹ ��L����M��S�Ug������G�&�s�,��p�x��^k�@ħe3��9�yy�#��T�4�R@Eg ݞ�ǳ��P���.��i	���$��$dFH~����s�Ң�������O����ƾ��:��0����,ZY�N��ܝ�f�p,v��]Z_�rT���
�~���?̤��F~�٣�H �����2g��bc������5���c�E�g#fL�3��6���PE->�r� �*0��3b��]����J.�����-���<-9��C�ogtg�C!1����+uoQ[̐&#�f·�B�0��j��� %�6��PǈcJS�t�ڇ.��g���U�Ote�/_0[L�YY���ba���λ����U^�_�Z=�w�!P�vB��GϨ�N�=�� h�k����퇀���,$��ܤ$p ������9b�5��k��i�a�ȑ��ܝg<!�;W�X�\P�࠸����K:a�`j���Dd�B�d�G�w@�ƶ	݈��f�����3���Q���Կ�˽��6:��V��@P�O��O�&%<��g��?{�����'�o͍�+u��}���S6e��
����n>EN]&���QŠL�9�I�YaU��75Ey��ϗ�����{�7��2��㓔��%���O��$���Г��	k&f�ӵ���Q��H��;u0�*/[���Zx�5"�J�G�\
��;lr��@����8u R�TR؀Ϛa ���Ѭl#��Ġ+�A�����8�8���1]:�CRb'^;%�$�W=?��mPJ!9MM;\\R"�m��x�tS�Ё���=��;���{Bq���M��!%�1*�n%b끹zyL�k�kr2�?"�����.��d�U���$��`�q��I�+a�w���.{Ѱc~�M���b�?5̧#Q��̾G�oke�C-:�X� 2Uo <�$��$z\�C�����D9C�J���X�AR92{�R����ѡ�9"�7	�H�'�8���T���I,�r�������:w�"���L/��q��s~�� �sv���D//���Ass����5g��JY�AZ���QU�/.yo�Z�w���&o}�.H��W�	��(�`��:j�84��
zh�������~�v���ڒk�kd¸!!R�n�|�����HVeb��6����᤯41���9Z�n��hzbj����ֵ��=�B��˓P�E�~wK2Hv�;K�2�Ν;����Y�L�*hp̺6�!�3��?����w6X	I:::�[.�R�rJ����[U�`�F(G�l�P)��p�v�zn��	�z0d�g[V���>hf���چ�;`����D�}����|�,���?L��y ���	�=� w���P#O��yQl!��Ri4���f3�n0���7�RZ����x׭j�$FVǖ�"���Ƹ.�%L�>@�_j���L�m���޸���<���_�b<�����m�������~�CW���o�o̴�x/ڒ8t�ژ��y�ڿ�YRR��^)���t�͑B2��z~S$d�ſ�IheL<��͗N��;G[|6��Y�8`~�E)Dxccc��`�����W� �aP����<u][s��%7 ��IW�k��t�� ʷˣ+mX�@)�X2����}�G
tX�����B�(@R,!N��7��9
�Sx),��
��
�����G���p\�re�-����ij )���^�w���3%$���� �{m��~∣��_e��Z�ּ��t����_�#u+(3Oz�6���r��M@RC�t��}�3 �k׀��}�o�)%�`7�{�f2�@B|Lb�N����+���d@L��u�J Z�����H8ܭ�}L@}��`y{��]ףj�u�Ha��w�����B�	�j���ڵ�Z�;�c��٦`��O���R.Z��D�E&ޖ�6�:�%��͜��1�_6)�n[�7�A��Q����t���I�.���?�}c�.����%'�^�-U`L�.���2\ ���um�m�][��j���|I<���)����У��v�u�F>�W�){A�{�X	 M���f4	bȹ�����v�'>���؍�� >k6�w>d�H5ǚ���z`̪�LR�[�uSyyy{�x>t6� ��4��tE����[u��х�,uEbm���D���а���.�I�y��iruz\*t���[gee]3<�����fg�X�����Ii�ZqS�P���O<���A䵁]F���lN���dm�V��1�����AT(� �W?���=V�̗���Lr���Y��&�3���~߫�R���]�֐'�i�f_. �L��9�1%k�����WE�)���umdWN|�!wz�C�B<F�f�4��y�ھ�~S�l9L2�J�&���Wa�RT�X+�Q2p�T��q�o<@;f�X��+�cR�C��C��" [ؗ�VF�@�)���.�h��$I�r0�*Ր�#ץ��m�I����]?�#]F���:e�2�>�G�,a������w*.�,�lVY?�yXl��I��A�r���*7��L�%����<�*JJ��:*-�2�5&��jdzU���jO����33����gö�$[i\@@DԪ�����a�zVo2�~C$P'yxhBڥ�|�e�$���g��K�z�g�xi���_ _�3�T����rg�jE�WPaT�N��%$%!G���O���J��贿�"�wK��nH$,j�W4-i�Xʋao7tS�ww����O��_n�\�~��R�=�������[~e:�Z� 
�	u�����?L<f��V�I� ��y�V�ؐl�ȥ�:r�z�J]Ʋ�?�V|h#.X�L�����*cf�@Ĝ5���z@@`��������$a�=�K��O����^d]еY%�,�!Ց��`��?�-���k�cÞ]�H�p��4Q�MM�6W����a5=Ыe���ސl&�lhmݔ��w�%[�p��u�)Ӣ��2V�H�c&�v����u��06p�����um���!���@�&�|�y�bZ���x����s�+�җ��
זoh�{��f����^�аu�n݃@�\p�/��%n�>z4}�n~h[��Ͼ�j��a'[���\�%75�Ng��юYO$�`ۏ�	��$��2�)�F� �����\Ⱥ6o���l�����Z���*Q�zSӪfn^> gt�j��5mh+�t�e��hր�rؗTu!ҳ�VX�ݺ����H�v_�C<(d����-I�z������Pb1�i�wD�w���k{���)
�HLJ�oooO�ص('p�����5������݇$CK�v���܀�`$���SO���zx�f�i��\G��Kg��*�e2���4_]�B�ބ��V �߉�xJr�Xj���1G¡��� �_ޟ6k-e�iw�?0A�1������V�<� X�27�.��,��5���^��i��{�R
�-ҳ�]��}�H\	�E���!�g$�����;R���)��E_�迄5��oJc�ϖ� gJjA6T4e�����wU��n�Og��ʾ��8
H.�k�%�Tx���������{i�_}\[PSG.8�ibe"1�2�f�L%��A����`)H��%T1H�S�1�!� �(�$r��J����#��B`����n��I���y�Ӟ������'��u/X�k�jbgQHA�/{�;�����?k��·kt��GQte��b�o�j��u���m���h��p�J�.ݰF7�n�=�+Dt-,z�����Գ�Q��ϋ��<B�M�'��0��t�9Y�[�' �F���r�ɿ=��V�����~¥B�r��"u��6����%�p���x�4[�0Mۄ����F�7����B�_��G�dx!���īZG&l�A>(�5�DB��� 0t?�\�ݬ�e�_c�' "�� ��f�B�;]L���ڜ!gr���9�]{j�R_8qHHHD&L�!��FV0lf��G��ܸ+P�)E������nvE/�w�v�f+?Y�9�Qs�$O�|8�i�Qx�m,�U�����ϗ%�;�������@����N'�Sͪ��&㈮z��7�	�?�S/��1��_L�4�|�L�:%���'�ʇ�m����������$�l�\��D���.)|Mܠ��C���َw �{�y���h@��'�ۯ,KV�W�ZW�������xR��~�1���� ��2`Z%@�kX��Sخ	�V�P	���:�޾�}w��9�ьA���Bp��	Ϧ ���Qg	�KsZ��T�\�V$�-����nQ�~,&wF�rJӻ�p�䋐ƐK��Xn�k>=k���7�UGWvT��{�3��BT�*'��}�؅�Sw�߽$>_�o7����������8b%ؽ��>�][]�z���2� Tu(
\ݖb�tZ�ݾx}Y���x�T��K��V'Gmu�@ݥ�{�Auʹ�_�<�3�9�!��p�a�t�V�)v~��W�������[u�C���[�T���j���!��NA��կ�>�w��Ĳe2{���Fظ���c���PP�����k�+�܃m����C_�7�a��v�Zss�;U[��N��S�)����`���HR#0S��;Qv��U��of��C�f�jS��q[o�3W�Z�O�A{��y0lPA�q���j�����9��ּ����Tl�`�GMx3)�"�	�L���DՆ�3�7��^�n	<�CUF��Ff����G��-�w�`A�Y� ���*�D�y6d�N?й6O�T�g���\�o?�QbS����.V@����Z�o>�����<z�ǣ��fs�Q�e��lAϗyr�F"-p�qUTA�T�;z6��!+��^E�٥"�U�x�	mIq� i��Is����.~��Ħ��`)��u���'d�d�H�|�git�Fbh���"��t�?���b`�	�A!��5�~Ĩx��|���f�L�Υ@%���P�aq�D�0�=eB���2���8������QSc����d��b'W=d�Z��x"#�y5���PK   ��X��g �  ��     jsons/user_defined.json�\ߏ�6�W�K������fs�[\��h���PE%B����N�+���H���5EY��;��ב�q��7�!��m��|�/������
u��t6�V��r��AZ ~r�)�K�/����W�rQ��*T������Y�����
o�n�/W��6��n���4��^�^�n~f��N+G%T�"��c)i퉫$����cy����[o���������<H���D�Z��$�2��
\�Lq�x���5�a9}�[�vk�f��k��Z\Vo׫�C_�k�Z�,��M3o��. (�:�}�eaQ�]D-�1F�e��7�a�B����j����2�7�[��~��G�h�
)�T���/��nN�����ޑ��H����$}���ԑ��~�;2h��}���������u�(4��������O��ɂ!�v����v�ѕ�fM�V˻�Z7;n�q�5�%��ݢՅ�oڿ��v
�!��>,?]/.��w_�ܲ�]sߴ0��¿6ͪ�};٭O���bS;�ެ�� ���իM��\.�M{�����b�� �F1��K�)�� 8�PKT�ӍG��",�����n�������������ǎ������O�	�����U��
�D]��!p�t��&��@t-y�Z�'��z�NĞGq�R�T��`]�H'����	n8�7Xa4J#6�!\@a���D�@�?,�06r �OfQ�h��-���$�
*�XQ`x��9�����.��3d�j�t�幵j*&�
���]��0UZ[j)�\�sϨ�QP���<F]�f�
��Z��3A\	@<���b-K,hujf��ve%*BKPDHV+#�_����X���Ô���E��1&/��9iy�=
�r�0l
\�l_�q5��/.�
����P���R���:�ۧ�sO���}��8�î,5��(%��`� ���Rf_f_f_f_f_f_f_f_f_f�8�r��-a>�'�����M�WO�x���5�S.n��QQVBRi�A�9b�Ě�,��KY��TT�z�Z͙'�V@��z�2��j�'v.���WB��d�{�))�7h.���gnJ�h�ݬ�Z�C�p�a<�A��2f��0&��0r��ePPhc�m
EA<�."\�#��(�Rf����`R6���T�9|&�-(nO@��^1��s�3�'�P��!��3���	3�+���f$�B.jp.(�b�1r�Rn�&B��!��匣
�����+Ӌ`��2�g�LF�a݋`��%)f�h��`h&.�T��"	�]p8�1�Ƀ+n�8{y%�!"I�����I	�L�a?�~���1:	��B|k��r��"�"�V�@�p����0�		U@L�9+�!s�Q��� ȓv��m0	��3���k��0ȓ���F)�(�&�J���	I�K��)ya���h�$5#�"o�
�5�֠MĠ!*9#�2o󒑘Pg(D��Ró���/��CI�V3�����&���E28JO��1�Sc�Y��&��tK���Y5�-}�:h�J�����%w1Q!����ǖ�f$�ȭ���$ӶU���I�HD�-��v&Ӆ�Xc��I�ds�PmѤ1]a�1����~&�1�J*D�'=&ud�D��$U��T��ĤA"Z�[�c<��8lIbFx4���	-0�bT)pu"�4�:��ќ�k��lh1fC
���~�c�#��X(������C%��+�q,�ne��ĺ�=Fk�1���̑�������ߕa��<�i&�Փ��M�WK�׫�|�nwZ�U��j��qo��$�����CU�S�[�7�(R�Za�/%)A���+��Pr�N���JQ,S�=���bԗH<�6!��:��#�P1���¹���'�1��9 ��Z�п�>N\z4@"��,s�����:�X��9�G��+zD?�"�
Zc���]?�"���5tL�	[-��mh1���4�g�h�������c._��6Y��tj����,F;e+�Q�݌�ZԞc$Dlci;�̀k#[Kp��X�W�ͥ�Ou�F��{ �����Έ~�EJ�G���R���`�G`@�d�
�=qO�HMFD��GAbe�~V#b��XF�q��8Zi�C���A���@��LǪ�}b#��p�2a���՘+�1F�/e#E��BmFb=~�m��~:��9���?V�>"A�cm��v���cm��vj"��=Z��]��E��y�	;'�Os�ɛ�ׯ�o_����Wo�B+���3�?jl ꝡ���K���B"B(C骠$�m5������ػ�+�F
~��l�Q��g@,hG�PׄU�'�Z��DU��ɧkQy�DR�B�51L�R*��e�N Pd�%c�3PHη��q�SF!a�I9�Ô�G����F���#��B�����<CNQ���!�}E�.�!���I}G'�hk��Y4_���E�`�]��h�#�R�y����9}2�B�4�eI�+�]sEJ鑺D������7YPź����ԃm?�Hz���]�K5���r$���KuO�R$����e�5Ly�.m�l �W�SF��~>v夙�f����������o�OL���5��.��<��paH�k&���!5�8���K]S�ik;fmr:hN�²�0�?���y���)ceYK���x��m�_R⃯�t���p>�BI�M��~�����"����m_�l;^�YG{@�i|U\�D+m
�k(�fz�����M"�纇 #
fԠ:������/�U�?�0Զٹ�c7r���0� \��~�ȉ�Ba��L�PT�~�ȡ�C�H�j�GX:W�ENU��5���d�uո~��`�~g��T?D�T��o-O�T���W�!@�0ZG% z%�\��b�k0��ƵD(�3���P���}�l�:���\� ��mb��n�@�0vp�i�tǀ�k�ػK�q׸戽���~�%��������F��GE��K��5��$уQ��]zg�P�jAR����5
dT�ā���]���I�G�w����$K�k�ػkHbyU<�r�e]Z�"�%v,��*q�ahۙ��ӈA&/�P�jT�D��:$ke�-����U"�ǚ&���c���a��"�?���R	;Ԟ�	zE$�!�)@ C��Ώˬ���-^�z��zI�B�DɈ�XVP����8QP;'P���'��9��	A�o�Ą��BYV����27]A�+]�nլ?oM�;�g��y8^�_דr���E��ೈ�7���z9	U�n���½��_�����R;����Ϧ����x�e������Gt7a]:����r����\w��o��4�b��s��Q0�Q���FEJ�Q���������`0�G�b�Y5a5�
�R�y�m�J�*���9-�* ��&0n1Ii���GӲ����������������������������������������������������������������������������������������������������������������������PK
   ��X�ji՗6  ��                  cirkitFile.jsonPK
   �sX��k��E  �E  /             �6  images/022bbf54-c303-4c74-b4b0-cecd35afa1b1.pngPK
   ��X���  �  /             �|  images/10ca8052-f8e9-4304-b468-4eebebade650.pngPK
   �sXUs?��B  0 /             3�  images/1e112c27-401d-49ee-8ccd-a7b22cee0ece.pngPK
   ��X����7  �  /             E� images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   �sX,�׳A}  7}  /             �� images/3d46b7b2-3c4d-4bbd-b0e2-e734cbc728a9.pngPK
   ��X�z��kW S� /             Wm images/65d233e5-7445-4b75-a6a5-2d8c2ad1af28.pngPK
   �sX��G��D [ /             � images/6e0c1376-732c-4f61-beca-ab02432631e3.pngPK
   ��X�1.:�  )  /             
 images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   �sX�@M��  2�  /             ") images/959826c8-9748-429e-bc6c-0234da684cdf.pngPK
   ��X�� �f  y�  /             -� images/96fabd4d-0b16-452b-94e2-688cfcbce531.pngPK
   �sX�X�޿� X /             W images/97f4dc10-5048-4749-8251-75563a783bed.pngPK
   ��X�&�}[  y`  /             c� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   ��X��g)�
  �
  /             -A images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.pngPK
   ��X�р0G3 �	 /             ]L images/cc0c8c86-b3f6-4855-b14e-2ffc61d63776.pngPK
   ��X�GDU7� �� /             � images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   ��X�|�	  	  /             uc images/e1d4e862-170d-4bac-8b1a-e4319ef50e6b.pngPK
   �sX���F�� % /             �l images/e299bea7-de73-4651-8213-9be9a85bbb4e.pngPK
   �sX�Rr5�  5 /             j images/ed2720bb-136d-4736-b5c1-9714f7ccc33b.pngPK
   ��X��g �  ��               � jsons/user_defined.jsonPK        �   